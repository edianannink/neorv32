-- #################################################################################################
-- # << NEORV32 - Main VHDL Package File (CPU and SoC) >>                                          #
-- # ********************************************************************************************* #
-- # BSD 3-Clause License                                                                          #
-- #                                                                                               #
-- # Copyright (c) 2023, Stephan Nolting. All rights reserved.                                     #
-- #                                                                                               #
-- # Redistribution and use in source and binary forms, with or without modification, are          #
-- # permitted provided that the following conditions are met:                                     #
-- #                                                                                               #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of        #
-- #    conditions and the following disclaimer.                                                   #
-- #                                                                                               #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of     #
-- #    conditions and the following disclaimer in the documentation and/or other materials        #
-- #    provided with the distribution.                                                            #
-- #                                                                                               #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to  #
-- #    endorse or promote products derived from this software without specific prior written      #
-- #    permission.                                                                                #
-- #                                                                                               #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS   #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF               #
-- # MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE    #
-- # COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     #
-- # EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE #
-- # GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED    #
-- # AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING     #
-- # NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED  #
-- # OF THE POSSIBILITY OF SUCH DAMAGE.                                                            #
-- # ********************************************************************************************* #
-- # The NEORV32 RISC-V Processor - https://github.com/stnolting/neorv32       (c) Stephan Nolting #
-- #################################################################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package neorv32_package is

-- ****************************************************************************************************************************
-- Architecture Configuration and Constants
-- ****************************************************************************************************************************

  -- Architecture Configuration -------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- max response time for processor-internal bus transactions --
  -- = cycles after which an *unacknowledged* internal bus access will timeout triggering a bus fault exception
  constant bus_timeout_c : natural := 15; -- default = 15

  -- instruction prefetch buffer depth --
  constant ipb_depth_c : natural := 2; -- hast to be a power of two, min 2, default 2

  -- instruction monitor: raise exception if multi-cycle operation times out --
  constant monitor_mc_tmo_c : natural := 9; -- = log2 of max execution cycles (default = 512 cycles)

  -- Architecture Constants -----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant hw_version_c : std_ulogic_vector(31 downto 0) := x"01090200"; -- hardware version
  constant archid_c     : natural := 19; -- official RISC-V architecture ID
  constant XLEN         : natural := 32; -- native data path width, do not change!

  -- Check if we're inside the Matrix -------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant is_simulation_c : boolean := false -- seems like we're on real hardware
-- pragma translate_off
-- synthesis translate_off
-- RTL_SYNTHESIS OFF
  or true -- this MIGHT be a simulation
-- RTL_SYNTHESIS ON
-- synthesis translate_on
-- pragma translate_on
  ;

-- ****************************************************************************************************************************
-- Processor Address Space Layout
-- ****************************************************************************************************************************

  -- Main Address Regions ---
  constant mem_imem_base_c : std_ulogic_vector(31 downto 0) := x"00000000"; -- IMEM size via generic
  constant mem_dmem_base_c : std_ulogic_vector(31 downto 0) := x"80000000"; -- DMEM size via generic
  constant mem_xip_base_c  : std_ulogic_vector(31 downto 0) := x"e0000000"; -- page (4MSBs) only!
  constant mem_xip_size_c  : natural := 256*1024*1024;
  constant mem_boot_base_c : std_ulogic_vector(31 downto 0) := x"ffffc000";
  constant mem_boot_size_c : natural := 8*1024;
  constant mem_io_base_c   : std_ulogic_vector(31 downto 0) := x"ffffe000";
  constant mem_io_size_c   : natural := 8*1024;

  -- Start of uncached memory access (256MB page / 4MSBs only) --
  constant uncached_begin_c  : std_ulogic_vector(31 downto 0) := x"f0000000";

  -- IO Address Map --
  constant iodev_size_c      : natural := 256; -- size of a single IO device (bytes)
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe000"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe100"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe200"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe300"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe400"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe500"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe600"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe700"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe800"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe900"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffea00"; -- reserved
  constant base_io_cfs_c     : std_ulogic_vector(31 downto 0) := x"ffffeb00";
  constant base_io_slink_c   : std_ulogic_vector(31 downto 0) := x"ffffec00";
  constant base_io_dma_c     : std_ulogic_vector(31 downto 0) := x"ffffed00";
  constant base_io_crc_c     : std_ulogic_vector(31 downto 0) := x"ffffee00";
  constant base_io_xip_c     : std_ulogic_vector(31 downto 0) := x"ffffef00";
  constant base_io_pwm_c     : std_ulogic_vector(31 downto 0) := x"fffff000";
  constant base_io_gptmr_c   : std_ulogic_vector(31 downto 0) := x"fffff100";
  constant base_io_onewire_c : std_ulogic_vector(31 downto 0) := x"fffff200";
  constant base_io_xirq_c    : std_ulogic_vector(31 downto 0) := x"fffff300";
  constant base_io_mtime_c   : std_ulogic_vector(31 downto 0) := x"fffff400";
  constant base_io_uart0_c   : std_ulogic_vector(31 downto 0) := x"fffff500";
  constant base_io_uart1_c   : std_ulogic_vector(31 downto 0) := x"fffff600";
  constant base_io_sdi_c     : std_ulogic_vector(31 downto 0) := x"fffff700";
  constant base_io_spi_c     : std_ulogic_vector(31 downto 0) := x"fffff800";
  constant base_io_twi_c     : std_ulogic_vector(31 downto 0) := x"fffff900";
  constant base_io_trng_c    : std_ulogic_vector(31 downto 0) := x"fffffa00";
  constant base_io_wdt_c     : std_ulogic_vector(31 downto 0) := x"fffffb00";
  constant base_io_gpio_c    : std_ulogic_vector(31 downto 0) := x"fffffc00";
  constant base_io_neoled_c  : std_ulogic_vector(31 downto 0) := x"fffffd00";
  constant base_io_sysinfo_c : std_ulogic_vector(31 downto 0) := x"fffffe00";
  constant base_io_dm_c      : std_ulogic_vector(31 downto 0) := x"ffffff00";

  -- On-Chip Debugger - Debug Module Entry Points (Code ROM) --
  constant dm_exc_entry_c  : std_ulogic_vector(31 downto 0) := x"ffffff00"; -- = base_io_dm_c + 0, exceptions entry point
  constant dm_park_entry_c : std_ulogic_vector(31 downto 0) := x"ffffff08"; -- = base_io_dm_c + 8, normal entry point

-- ****************************************************************************************************************************
-- SoC Definitions
-- ****************************************************************************************************************************

  -- SoC Clock Select -----------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant clk_div2_c    : natural := 0;
  constant clk_div4_c    : natural := 1;
  constant clk_div8_c    : natural := 2;
  constant clk_div64_c   : natural := 3;
  constant clk_div128_c  : natural := 4;
  constant clk_div1024_c : natural := 5;
  constant clk_div2048_c : natural := 6;
  constant clk_div4096_c : natural := 7;

  -- Internal Memory Types ------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  type mem32_t is array (natural range <>) of std_ulogic_vector(31 downto 0); -- memory with 32-bit entries
  type mem16_t is array (natural range <>) of std_ulogic_vector(15 downto 0); -- memory with 16-bit entries
  type mem8_t  is array (natural range <>) of std_ulogic_vector(07 downto 0); -- memory with 8-bit entries
  
  type mem15_t  is array (natural range <>) of std_ulogic_vector(14 downto 0); -- memory with 15-bit entries
  type mem13_t  is array (natural range <>) of std_ulogic_vector(12 downto 0); -- memory with 13-bit entries

  -- Internal Bus Interface -----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- bus request --
  type bus_req_t is record
    addr : std_ulogic_vector(31 downto 0); -- access address
    data : std_ulogic_vector(31 downto 0); -- write data
    ben  : std_ulogic_vector(03 downto 0); -- byte enable
    stb  : std_ulogic; -- request strobe (single-shot)
    rw   : std_ulogic; -- 0=read, 1=write
    src  : std_ulogic; -- access source (1=instruction fetch, 0=data access)
    priv : std_ulogic; -- set if privileged (machine-mode) access
    rvso : std_ulogic; -- set if reservation set operation (atomic LR/SC)
  end record;

  -- bus response --
  type bus_rsp_t is record
    data : std_ulogic_vector(31 downto 0); -- read data
    ack  : std_ulogic; -- access acknowledge (single-shot)
    err  : std_ulogic; -- access error (single-shot)
  end record;

  -- source (request) termination --
  constant req_terminate_c : bus_req_t := (
    addr => (others => '0'),
    data => (others => '0'),
    ben  => (others => '0'),
    stb  => '0',
    rw   => '0',
    src  => '0',
    priv => '0',
    rvso => '0'
  );

  -- endpoint (response) termination --
  constant rsp_terminate_c : bus_rsp_t := (
    data => (others => '0'),
    ack  => '0',
    err  => '0'
  );

  -- Debug Module Interface -----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- request --
  type dmi_req_t is record
    addr : std_ulogic_vector(06 downto 0);
    op   : std_ulogic_vector(01 downto 0);
    data : std_ulogic_vector(31 downto 0);
  end record;

  -- request operation --
  constant dmi_req_nop_c : std_ulogic_vector(1 downto 0) := "00"; -- no operation
  constant dmi_req_rd_c  : std_ulogic_vector(1 downto 0) := "01"; -- read access
  constant dmi_req_wr_c  : std_ulogic_vector(1 downto 0) := "10"; -- write access

  -- response --
  type dmi_rsp_t is record
    data : std_ulogic_vector(31 downto 0);
    ack  : std_ulogic;
  end record;

-- ****************************************************************************************************************************
-- RISC-V ISA Definitions
-- ****************************************************************************************************************************

  -- RISC-V 32-Bit Instruction Word Layout --------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant instr_opcode_lsb_c  : natural :=  0; -- opcode bit 0
  constant instr_opcode_msb_c  : natural :=  6; -- opcode bit 6
  constant instr_rd_lsb_c      : natural :=  7; -- destination register address bit 0
  constant instr_rd_msb_c      : natural := 11; -- destination register address bit 4
  constant instr_funct3_lsb_c  : natural := 12; -- funct3 bit 0
  constant instr_funct3_msb_c  : natural := 14; -- funct3 bit 2
  constant instr_rs1_lsb_c     : natural := 15; -- source register 1 address bit 0
  constant instr_rs1_msb_c     : natural := 19; -- source register 1 address bit 4
  constant instr_rs2_lsb_c     : natural := 20; -- source register 2 address bit 0
  constant instr_rs2_msb_c     : natural := 24; -- source register 2 address bit 4
  constant instr_rs3_lsb_c     : natural := 27; -- source register 3 address bit 0
  constant instr_rs3_msb_c     : natural := 31; -- source register 3 address bit 4
  constant instr_funct7_lsb_c  : natural := 25; -- funct7 bit 0
  constant instr_funct7_msb_c  : natural := 31; -- funct7 bit 6
  constant instr_funct12_lsb_c : natural := 20; -- funct12 bit 0
  constant instr_funct12_msb_c : natural := 31; -- funct12 bit 11
  constant instr_imm12_lsb_c   : natural := 20; -- immediate12 bit 0
  constant instr_imm12_msb_c   : natural := 31; -- immediate12 bit 11
  constant instr_imm20_lsb_c   : natural := 12; -- immediate20 bit 0
  constant instr_imm20_msb_c   : natural := 31; -- immediate20 bit 21
  constant instr_funct5_lsb_c  : natural := 27; -- funct5 select bit 0
  constant instr_funct5_msb_c  : natural := 31; -- funct5 select bit 4

  -- RISC-V Opcodes -------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- alu --
  constant opcode_alui_c   : std_ulogic_vector(6 downto 0) := "0010011"; -- ALU operation with immediate
  constant opcode_alu_c    : std_ulogic_vector(6 downto 0) := "0110011"; -- ALU operation
  constant opcode_lui_c    : std_ulogic_vector(6 downto 0) := "0110111"; -- load upper immediate
  constant opcode_auipc_c  : std_ulogic_vector(6 downto 0) := "0010111"; -- add upper immediate to PC
  -- control flow --
  constant opcode_jal_c    : std_ulogic_vector(6 downto 0) := "1101111"; -- jump and link
  constant opcode_jalr_c   : std_ulogic_vector(6 downto 0) := "1100111"; -- jump and link with register
  constant opcode_branch_c : std_ulogic_vector(6 downto 0) := "1100011"; -- branch
  -- memory access --
  constant opcode_load_c   : std_ulogic_vector(6 downto 0) := "0000011"; -- load
  constant opcode_store_c  : std_ulogic_vector(6 downto 0) := "0100011"; -- store
  constant opcode_amo_c    : std_ulogic_vector(6 downto 0) := "0101111"; -- atomic memory access
  constant opcode_fence_c  : std_ulogic_vector(6 downto 0) := "0001111"; -- fence / fence.i
  -- system/csr --
  constant opcode_system_c : std_ulogic_vector(6 downto 0) := "1110011"; -- system/csr access
  -- floating point operations --
  constant opcode_fop_c    : std_ulogic_vector(6 downto 0) := "1010011"; -- dual/single operand instruction
  -- official custom RISC-V opcodes - free for custom instructions --
  constant opcode_cust0_c  : std_ulogic_vector(6 downto 0) := "0001011"; -- custom-0
  constant opcode_cust1_c  : std_ulogic_vector(6 downto 0) := "0101011"; -- custom-1
  constant opcode_cust2_c  : std_ulogic_vector(6 downto 0) := "1011011"; -- custom-2
  constant opcode_cust3_c  : std_ulogic_vector(6 downto 0) := "1111011"; -- custom-3

  -- RISC-V Funct3 --------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- control flow --
  constant funct3_beq_c    : std_ulogic_vector(2 downto 0) := "000"; -- branch if equal
  constant funct3_bne_c    : std_ulogic_vector(2 downto 0) := "001"; -- branch if not equal
  constant funct3_blt_c    : std_ulogic_vector(2 downto 0) := "100"; -- branch if less than
  constant funct3_bge_c    : std_ulogic_vector(2 downto 0) := "101"; -- branch if greater than or equal
  constant funct3_bltu_c   : std_ulogic_vector(2 downto 0) := "110"; -- branch if less than (unsigned)
  constant funct3_bgeu_c   : std_ulogic_vector(2 downto 0) := "111"; -- branch if greater than or equal (unsigned)
  -- memory access --
  constant funct3_lb_c     : std_ulogic_vector(2 downto 0) := "000"; -- load byte (signed)
  constant funct3_lh_c     : std_ulogic_vector(2 downto 0) := "001"; -- load half word (signed)
  constant funct3_lw_c     : std_ulogic_vector(2 downto 0) := "010"; -- load word (signed)
  constant funct3_lbu_c    : std_ulogic_vector(2 downto 0) := "100"; -- load byte (unsigned)
  constant funct3_lhu_c    : std_ulogic_vector(2 downto 0) := "101"; -- load half word (unsigned)
  constant funct3_lwu_c    : std_ulogic_vector(2 downto 0) := "110"; -- load word (unsigned)
  constant funct3_sb_c     : std_ulogic_vector(2 downto 0) := "000"; -- store byte
  constant funct3_sh_c     : std_ulogic_vector(2 downto 0) := "001"; -- store half word
  constant funct3_sw_c     : std_ulogic_vector(2 downto 0) := "010"; -- store word
  -- alu --
  constant funct3_subadd_c : std_ulogic_vector(2 downto 0) := "000"; -- sub/add via funct7
  constant funct3_sll_c    : std_ulogic_vector(2 downto 0) := "001"; -- shift logical left
  constant funct3_slt_c    : std_ulogic_vector(2 downto 0) := "010"; -- set on less
  constant funct3_sltu_c   : std_ulogic_vector(2 downto 0) := "011"; -- set on less unsigned
  constant funct3_xor_c    : std_ulogic_vector(2 downto 0) := "100"; -- xor
  constant funct3_sr_c     : std_ulogic_vector(2 downto 0) := "101"; -- shift right via funct7
  constant funct3_or_c     : std_ulogic_vector(2 downto 0) := "110"; -- or
  constant funct3_and_c    : std_ulogic_vector(2 downto 0) := "111"; -- and
  -- system/csr --
  constant funct3_env_c    : std_ulogic_vector(2 downto 0) := "000"; -- ecall, ebreak, mret, wfi, ...
  constant funct3_csrrw_c  : std_ulogic_vector(2 downto 0) := "001"; -- csr r/w
  constant funct3_csrrs_c  : std_ulogic_vector(2 downto 0) := "010"; -- csr read & set
  constant funct3_csrrc_c  : std_ulogic_vector(2 downto 0) := "011"; -- csr read & clear
  constant funct3_csril_c  : std_ulogic_vector(2 downto 0) := "100"; -- undefined/illegal csr command
  constant funct3_csrrwi_c : std_ulogic_vector(2 downto 0) := "101"; -- csr r/w immediate
  constant funct3_csrrsi_c : std_ulogic_vector(2 downto 0) := "110"; -- csr read & set immediate
  constant funct3_csrrci_c : std_ulogic_vector(2 downto 0) := "111"; -- csr read & clear immediate
  -- fence --
  constant funct3_fence_c  : std_ulogic_vector(2 downto 0) := "000"; -- fence - order IO/memory access
  constant funct3_fencei_c : std_ulogic_vector(2 downto 0) := "001"; -- fence.i - instruction stream sync

  -- RISC-V Funct12 - SYSTEM ----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant funct12_ecall_c  : std_ulogic_vector(11 downto 0) := x"000"; -- ecall
  constant funct12_ebreak_c : std_ulogic_vector(11 downto 0) := x"001"; -- ebreak
  constant funct12_wfi_c    : std_ulogic_vector(11 downto 0) := x"105"; -- wfi
  constant funct12_mret_c   : std_ulogic_vector(11 downto 0) := x"302"; -- mret
  constant funct12_dret_c   : std_ulogic_vector(11 downto 0) := x"7b2"; -- dret

  -- RISC-V Floating-Point Stuff ------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant float_single_c : std_ulogic_vector(1 downto 0) := "00"; -- single-precision (32-bit)
--constant float_double_c : std_ulogic_vector(1 downto 0) := "01"; -- double-precision (64-bit)
--constant float_half_c   : std_ulogic_vector(1 downto 0) := "10"; -- half-precision (16-bit)
--constant float_quad_c   : std_ulogic_vector(1 downto 0) := "11"; -- quad-precision (128-bit)

  -- number class flags --
  constant fp_class_neg_inf_c    : natural := 0; -- negative infinity
  constant fp_class_neg_norm_c   : natural := 1; -- negative normal number
  constant fp_class_neg_denorm_c : natural := 2; -- negative subnormal number
  constant fp_class_neg_zero_c   : natural := 3; -- negative zero
  constant fp_class_pos_zero_c   : natural := 4; -- positive zero
  constant fp_class_pos_denorm_c : natural := 5; -- positive subnormal number
  constant fp_class_pos_norm_c   : natural := 6; -- positive normal number
  constant fp_class_pos_inf_c    : natural := 7; -- positive infinity
  constant fp_class_snan_c       : natural := 8; -- signaling NaN (sNaN)
  constant fp_class_qnan_c       : natural := 9; -- quiet NaN (qNaN)

  -- exception flags --
  constant fp_exc_nx_c : natural := 0; -- inexact
  constant fp_exc_uf_c : natural := 1; -- underflow
  constant fp_exc_of_c : natural := 2; -- overflow
  constant fp_exc_dz_c : natural := 3; -- division by zero
  constant fp_exc_nv_c : natural := 4; -- invalid operation

  -- special values (single-precision) --
  constant fp_single_qnan_c     : std_ulogic_vector(31 downto 0) := x"7fc00000"; -- quiet NaN
  constant fp_single_snan_c     : std_ulogic_vector(31 downto 0) := x"7fa00000"; -- signaling NaN
  constant fp_single_pos_inf_c  : std_ulogic_vector(31 downto 0) := x"7f800000"; -- positive infinity
  constant fp_single_neg_inf_c  : std_ulogic_vector(31 downto 0) := x"ff800000"; -- negative infinity
  constant fp_single_pos_zero_c : std_ulogic_vector(31 downto 0) := x"00000000"; -- positive zero
  constant fp_single_neg_zero_c : std_ulogic_vector(31 downto 0) := x"80000000"; -- negative zero

  -- RISC-V CSRs ----------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- user floating-point CSRs --
  constant csr_fflags_c         : std_ulogic_vector(11 downto 0) := x"001";
  constant csr_frm_c            : std_ulogic_vector(11 downto 0) := x"002";
  constant csr_fcsr_c           : std_ulogic_vector(11 downto 0) := x"003";
  -- machine trap setup --
  constant csr_mstatus_c        : std_ulogic_vector(11 downto 0) := x"300";
  constant csr_misa_c           : std_ulogic_vector(11 downto 0) := x"301";
  constant csr_mie_c            : std_ulogic_vector(11 downto 0) := x"304";
  constant csr_mtvec_c          : std_ulogic_vector(11 downto 0) := x"305";
  constant csr_mcounteren_c     : std_ulogic_vector(11 downto 0) := x"306";
  constant csr_mstatush_c       : std_ulogic_vector(11 downto 0) := x"310";
  -- machine configuration --
  constant csr_menvcfg_c        : std_ulogic_vector(11 downto 0) := x"30a";
  constant csr_menvcfgh_c       : std_ulogic_vector(11 downto 0) := x"31a";
  -- machine counter setup --
  constant csr_mcountinhibit_c  : std_ulogic_vector(11 downto 0) := x"320";
  constant csr_mcyclecfg_c      : std_ulogic_vector(11 downto 0) := x"321";
  constant csr_minstretcfg_c    : std_ulogic_vector(11 downto 0) := x"322";
  constant csr_mhpmevent3_c     : std_ulogic_vector(11 downto 0) := x"323";
  constant csr_mhpmevent4_c     : std_ulogic_vector(11 downto 0) := x"324";
  constant csr_mhpmevent5_c     : std_ulogic_vector(11 downto 0) := x"325";
  constant csr_mhpmevent6_c     : std_ulogic_vector(11 downto 0) := x"326";
  constant csr_mhpmevent7_c     : std_ulogic_vector(11 downto 0) := x"327";
  constant csr_mhpmevent8_c     : std_ulogic_vector(11 downto 0) := x"328";
  constant csr_mhpmevent9_c     : std_ulogic_vector(11 downto 0) := x"329";
  constant csr_mhpmevent10_c    : std_ulogic_vector(11 downto 0) := x"32a";
  constant csr_mhpmevent11_c    : std_ulogic_vector(11 downto 0) := x"32b";
  constant csr_mhpmevent12_c    : std_ulogic_vector(11 downto 0) := x"32c";
  constant csr_mhpmevent13_c    : std_ulogic_vector(11 downto 0) := x"32d";
  constant csr_mhpmevent14_c    : std_ulogic_vector(11 downto 0) := x"32e";
  constant csr_mhpmevent15_c    : std_ulogic_vector(11 downto 0) := x"32f";
  -- machine trap handling --
  constant csr_mscratch_c       : std_ulogic_vector(11 downto 0) := x"340";
  constant csr_mepc_c           : std_ulogic_vector(11 downto 0) := x"341";
  constant csr_mcause_c         : std_ulogic_vector(11 downto 0) := x"342";
  constant csr_mtval_c          : std_ulogic_vector(11 downto 0) := x"343";
  constant csr_mip_c            : std_ulogic_vector(11 downto 0) := x"344";
  constant csr_mtinst_c         : std_ulogic_vector(11 downto 0) := x"34a";
  -- physical memory protection - configuration --
  constant csr_pmpcfg0_c        : std_ulogic_vector(11 downto 0) := x"3a0";
  constant csr_pmpcfg1_c        : std_ulogic_vector(11 downto 0) := x"3a1";
  constant csr_pmpcfg2_c        : std_ulogic_vector(11 downto 0) := x"3a2";
  constant csr_pmpcfg3_c        : std_ulogic_vector(11 downto 0) := x"3a3";
  -- physical memory protection - address --
  constant csr_pmpaddr0_c       : std_ulogic_vector(11 downto 0) := x"3b0";
  constant csr_pmpaddr1_c       : std_ulogic_vector(11 downto 0) := x"3b1";
  constant csr_pmpaddr2_c       : std_ulogic_vector(11 downto 0) := x"3b2";
  constant csr_pmpaddr3_c       : std_ulogic_vector(11 downto 0) := x"3b3";
  constant csr_pmpaddr4_c       : std_ulogic_vector(11 downto 0) := x"3b4";
  constant csr_pmpaddr5_c       : std_ulogic_vector(11 downto 0) := x"3b5";
  constant csr_pmpaddr6_c       : std_ulogic_vector(11 downto 0) := x"3b6";
  constant csr_pmpaddr7_c       : std_ulogic_vector(11 downto 0) := x"3b7";
  constant csr_pmpaddr8_c       : std_ulogic_vector(11 downto 0) := x"3b8";
  constant csr_pmpaddr9_c       : std_ulogic_vector(11 downto 0) := x"3b9";
  constant csr_pmpaddr10_c      : std_ulogic_vector(11 downto 0) := x"3ba";
  constant csr_pmpaddr11_c      : std_ulogic_vector(11 downto 0) := x"3bb";
  constant csr_pmpaddr12_c      : std_ulogic_vector(11 downto 0) := x"3bc";
  constant csr_pmpaddr13_c      : std_ulogic_vector(11 downto 0) := x"3bd";
  constant csr_pmpaddr14_c      : std_ulogic_vector(11 downto 0) := x"3be";
  constant csr_pmpaddr15_c      : std_ulogic_vector(11 downto 0) := x"3bf";
  -- machine counter setup - continued --
  constant csr_mcyclecfgh_c     : std_ulogic_vector(11 downto 0) := x"721";
  constant csr_minstretcfgh_c   : std_ulogic_vector(11 downto 0) := x"722";
  -- trigger module registers --
  constant csr_tselect_c        : std_ulogic_vector(11 downto 0) := x"7a0";
  constant csr_tdata1_c         : std_ulogic_vector(11 downto 0) := x"7a1";
  constant csr_tdata2_c         : std_ulogic_vector(11 downto 0) := x"7a2";
  constant csr_tinfo_c          : std_ulogic_vector(11 downto 0) := x"7a4";
  -- debug mode registers --
  constant csr_dcsr_c           : std_ulogic_vector(11 downto 0) := x"7b0";
  constant csr_dpc_c            : std_ulogic_vector(11 downto 0) := x"7b1";
  constant csr_dscratch0_c      : std_ulogic_vector(11 downto 0) := x"7b2";
  -- NEORV32-specific (user-mode) registers --
  constant csr_cfureg0_c        : std_ulogic_vector(11 downto 0) := x"800";
  constant csr_cfureg1_c        : std_ulogic_vector(11 downto 0) := x"801";
  constant csr_cfureg2_c        : std_ulogic_vector(11 downto 0) := x"802";
  constant csr_cfureg3_c        : std_ulogic_vector(11 downto 0) := x"803";
  -- machine counters/timers --
  constant csr_mcycle_c         : std_ulogic_vector(11 downto 0) := x"b00";
--constant csr_mtime_c          : std_ulogic_vector(11 downto 0) := x"b01";
  constant csr_minstret_c       : std_ulogic_vector(11 downto 0) := x"b02";
  constant csr_mhpmcounter3_c   : std_ulogic_vector(11 downto 0) := x"b03";
  constant csr_mhpmcounter4_c   : std_ulogic_vector(11 downto 0) := x"b04";
  constant csr_mhpmcounter5_c   : std_ulogic_vector(11 downto 0) := x"b05";
  constant csr_mhpmcounter6_c   : std_ulogic_vector(11 downto 0) := x"b06";
  constant csr_mhpmcounter7_c   : std_ulogic_vector(11 downto 0) := x"b07";
  constant csr_mhpmcounter8_c   : std_ulogic_vector(11 downto 0) := x"b08";
  constant csr_mhpmcounter9_c   : std_ulogic_vector(11 downto 0) := x"b09";
  constant csr_mhpmcounter10_c  : std_ulogic_vector(11 downto 0) := x"b0a";
  constant csr_mhpmcounter11_c  : std_ulogic_vector(11 downto 0) := x"b0b";
  constant csr_mhpmcounter12_c  : std_ulogic_vector(11 downto 0) := x"b0c";
  constant csr_mhpmcounter13_c  : std_ulogic_vector(11 downto 0) := x"b0d";
  constant csr_mhpmcounter14_c  : std_ulogic_vector(11 downto 0) := x"b0e";
  constant csr_mhpmcounter15_c  : std_ulogic_vector(11 downto 0) := x"b0f";
  --
  constant csr_mcycleh_c        : std_ulogic_vector(11 downto 0) := x"b80";
--constant csr_mtimeh_c         : std_ulogic_vector(11 downto 0) := x"b81";
  constant csr_minstreth_c      : std_ulogic_vector(11 downto 0) := x"b82";
  constant csr_mhpmcounter3h_c  : std_ulogic_vector(11 downto 0) := x"b83";
  constant csr_mhpmcounter4h_c  : std_ulogic_vector(11 downto 0) := x"b84";
  constant csr_mhpmcounter5h_c  : std_ulogic_vector(11 downto 0) := x"b85";
  constant csr_mhpmcounter6h_c  : std_ulogic_vector(11 downto 0) := x"b86";
  constant csr_mhpmcounter7h_c  : std_ulogic_vector(11 downto 0) := x"b87";
  constant csr_mhpmcounter8h_c  : std_ulogic_vector(11 downto 0) := x"b88";
  constant csr_mhpmcounter9h_c  : std_ulogic_vector(11 downto 0) := x"b89";
  constant csr_mhpmcounter10h_c : std_ulogic_vector(11 downto 0) := x"b8a";
  constant csr_mhpmcounter11h_c : std_ulogic_vector(11 downto 0) := x"b8b";
  constant csr_mhpmcounter12h_c : std_ulogic_vector(11 downto 0) := x"b8c";
  constant csr_mhpmcounter13h_c : std_ulogic_vector(11 downto 0) := x"b8d";
  constant csr_mhpmcounter14h_c : std_ulogic_vector(11 downto 0) := x"b8e";
  constant csr_mhpmcounter15h_c : std_ulogic_vector(11 downto 0) := x"b8f";
  -- user counters/timers --
  constant csr_cycle_c          : std_ulogic_vector(11 downto 0) := x"c00";
  constant csr_time_c           : std_ulogic_vector(11 downto 0) := x"c01";
  constant csr_instret_c        : std_ulogic_vector(11 downto 0) := x"c02";
  constant csr_hpmcounter3_c    : std_ulogic_vector(11 downto 0) := x"c03";
  constant csr_hpmcounter4_c    : std_ulogic_vector(11 downto 0) := x"c04";
  constant csr_hpmcounter5_c    : std_ulogic_vector(11 downto 0) := x"c05";
  constant csr_hpmcounter6_c    : std_ulogic_vector(11 downto 0) := x"c06";
  constant csr_hpmcounter7_c    : std_ulogic_vector(11 downto 0) := x"c07";
  constant csr_hpmcounter8_c    : std_ulogic_vector(11 downto 0) := x"c08";
  constant csr_hpmcounter9_c    : std_ulogic_vector(11 downto 0) := x"c09";
  constant csr_hpmcounter10_c   : std_ulogic_vector(11 downto 0) := x"c0a";
  constant csr_hpmcounter11_c   : std_ulogic_vector(11 downto 0) := x"c0b";
  constant csr_hpmcounter12_c   : std_ulogic_vector(11 downto 0) := x"c0c";
  constant csr_hpmcounter13_c   : std_ulogic_vector(11 downto 0) := x"c0d";
  constant csr_hpmcounter14_c   : std_ulogic_vector(11 downto 0) := x"c0e";
  constant csr_hpmcounter15_c   : std_ulogic_vector(11 downto 0) := x"c0f";
  --
  constant csr_cycleh_c         : std_ulogic_vector(11 downto 0) := x"c80";
  constant csr_timeh_c          : std_ulogic_vector(11 downto 0) := x"c81";
  constant csr_instreth_c       : std_ulogic_vector(11 downto 0) := x"c82";
  constant csr_hpmcounter3h_c   : std_ulogic_vector(11 downto 0) := x"c83";
  constant csr_hpmcounter4h_c   : std_ulogic_vector(11 downto 0) := x"c84";
  constant csr_hpmcounter5h_c   : std_ulogic_vector(11 downto 0) := x"c85";
  constant csr_hpmcounter6h_c   : std_ulogic_vector(11 downto 0) := x"c86";
  constant csr_hpmcounter7h_c   : std_ulogic_vector(11 downto 0) := x"c87";
  constant csr_hpmcounter8h_c   : std_ulogic_vector(11 downto 0) := x"c88";
  constant csr_hpmcounter9h_c   : std_ulogic_vector(11 downto 0) := x"c89";
  constant csr_hpmcounter10h_c  : std_ulogic_vector(11 downto 0) := x"c8a";
  constant csr_hpmcounter11h_c  : std_ulogic_vector(11 downto 0) := x"c8b";
  constant csr_hpmcounter12h_c  : std_ulogic_vector(11 downto 0) := x"c8c";
  constant csr_hpmcounter13h_c  : std_ulogic_vector(11 downto 0) := x"c8d";
  constant csr_hpmcounter14h_c  : std_ulogic_vector(11 downto 0) := x"c8e";
  constant csr_hpmcounter15h_c  : std_ulogic_vector(11 downto 0) := x"c8f";
  -- machine information registers --
  constant csr_mvendorid_c      : std_ulogic_vector(11 downto 0) := x"f11";
  constant csr_marchid_c        : std_ulogic_vector(11 downto 0) := x"f12";
  constant csr_mimpid_c         : std_ulogic_vector(11 downto 0) := x"f13";
  constant csr_mhartid_c        : std_ulogic_vector(11 downto 0) := x"f14";
  constant csr_mconfigptr_c     : std_ulogic_vector(11 downto 0) := x"f15";
  -- NEORV32-specific (machine-mode) registers --
  constant csr_mxisa_c          : std_ulogic_vector(11 downto 0) := x"fc0";

-- ****************************************************************************************************************************
-- CPU Control
-- ****************************************************************************************************************************

  -- Main CPU Control Bus -------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  type ctrl_bus_t is record
    -- register file --
    rf_wb_en     : std_ulogic; -- write back enable
    rf_rs1       : std_ulogic_vector(04 downto 0); -- source register 1 address
    rf_rs2       : std_ulogic_vector(04 downto 0); -- source register 2 address
    rf_rs3       : std_ulogic_vector(04 downto 0); -- source register 3 address
    rf_rd        : std_ulogic_vector(04 downto 0); -- destination register address
    rf_mux       : std_ulogic_vector(01 downto 0); -- input source select
    rf_zero_we   : std_ulogic;                     -- allow/force write access to x0
    -- alu --
    alu_op       : std_ulogic_vector(02 downto 0); -- ALU operation select
    alu_opa_mux  : std_ulogic;                     -- operand A select (0=rs1, 1=PC)
    alu_opb_mux  : std_ulogic;                     -- operand B select (0=rs2, 1=IMM)
    alu_unsigned : std_ulogic;                     -- is unsigned ALU operation
    alu_cp_trig  : std_ulogic_vector(04 downto 0); -- co-processor trigger (one-hot)
    -- load/store unit --
    lsu_req      : std_ulogic;                     -- trigger memory access request
    lsu_rw       : std_ulogic;                     -- 0: read access, 1: write access
    lsu_mo_we    : std_ulogic;                     -- memory address and data output register write enable
    lsu_fence    : std_ulogic;                     -- fence operation
    lsu_fencei   : std_ulogic;                     -- fence.i operation
    lsu_priv     : std_ulogic;                     -- effective privilege level for load/store
    -- instruction word --
    ir_funct3    : std_ulogic_vector(02 downto 0); -- funct3 bit field
    ir_funct12   : std_ulogic_vector(11 downto 0); -- funct12 bit field
    ir_opcode    : std_ulogic_vector(06 downto 0); -- opcode bit field
    -- cpu status --
    cpu_priv     : std_ulogic;                     -- effective privilege mode
    cpu_sleep    : std_ulogic;                     -- set when CPU is in sleep mode
    cpu_trap     : std_ulogic;                     -- set when CPU is entering trap exec
    cpu_debug    : std_ulogic;                     -- set when CPU is in debug mode
  end record;

  -- control bus reset initializer --
  constant ctrl_bus_zero_c : ctrl_bus_t := (
    rf_wb_en     => '0',
    rf_rs1       => (others => '0'),
    rf_rs2       => (others => '0'),
    rf_rs3       => (others => '0'),
    rf_rd        => (others => '0'),
    rf_mux       => (others => '0'),
    rf_zero_we   => '0',
    alu_op       => (others => '0'),
    alu_opa_mux  => '0',
    alu_opb_mux  => '0',
    alu_unsigned => '0',
    alu_cp_trig  => (others => '0'),
    lsu_req      => '0',
    lsu_rw       => '0',
    lsu_mo_we    => '0',
    lsu_fence    => '0',
    lsu_fencei   => '0',
    lsu_priv     => '0',
    ir_funct3    => (others => '0'),
    ir_funct12   => (others => '0'),
    ir_opcode    => (others => '0'),
    cpu_priv     => '0',
    cpu_sleep    => '0',
    cpu_trap     => '0',
    cpu_debug    => '0'
  );

  -- Comparator Bus -------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant cmp_equal_c : natural := 0;
  constant cmp_less_c  : natural := 1; -- for signed and unsigned comparisons

  -- CPU Co-Processor IDs -------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant cp_sel_shifter_c  : natural := 0; -- CP0: shift operations (base ISA)
  constant cp_sel_muldiv_c   : natural := 1; -- CP1: multiplication/division operations ('M' extensions)
  constant cp_sel_bitmanip_c : natural := 2; -- CP2: bit manipulation ('B' extensions)
  constant cp_sel_fpu_c      : natural := 3; -- CP3: floating-point unit ('Zfinx' extension)
  constant cp_sel_cfu_c      : natural := 4; -- CP4: custom instructions CFU ('Zxcfu' extension)

  -- ALU Function Codes [DO NOT CHANGE ENCODING!] -------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant alu_op_add_c  : std_ulogic_vector(2 downto 0) := "000"; -- result <= A + B
  constant alu_op_sub_c  : std_ulogic_vector(2 downto 0) := "001"; -- result <= A - B
  constant alu_op_cp_c   : std_ulogic_vector(2 downto 0) := "010"; -- result <= ALU co-processor
  constant alu_op_slt_c  : std_ulogic_vector(2 downto 0) := "011"; -- result <= A < B
  constant alu_op_movb_c : std_ulogic_vector(2 downto 0) := "100"; -- result <= B
  constant alu_op_xor_c  : std_ulogic_vector(2 downto 0) := "101"; -- result <= A xor B
  constant alu_op_or_c   : std_ulogic_vector(2 downto 0) := "110"; -- result <= A or B
  constant alu_op_and_c  : std_ulogic_vector(2 downto 0) := "111"; -- result <= A and B

  -- Register File Input Select -------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant rf_mux_alu_c : std_ulogic_vector(1 downto 0) := "00"; -- register file <= alu result
  constant rf_mux_mem_c : std_ulogic_vector(1 downto 0) := "01"; -- register file <= memory read data
  constant rf_mux_csr_c : std_ulogic_vector(1 downto 0) := "10"; -- register file <= CSR read data
  constant rf_mux_ret_c : std_ulogic_vector(1 downto 0) := "11"; -- register file <= link-PC (return address)

  -- Trap ID Codes --------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- MSB:   1 = interrupt, 0 = sync. exception
  -- MSB-1: 1 = entry to debug mode, 0 = normal trapping
  -- RISC-V compliant synchronous exceptions --
  constant trap_ima_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00000"; -- 0: instruction misaligned
  constant trap_iaf_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00001"; -- 1: instruction access fault
  constant trap_iil_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00010"; -- 2: illegal instruction
  constant trap_brk_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00011"; -- 3: breakpoint
  constant trap_lma_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00100"; -- 4: load address misaligned
  constant trap_laf_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00101"; -- 5: load access fault
  constant trap_sma_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00110"; -- 6: store address misaligned
  constant trap_saf_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00111"; -- 7: store access fault
  constant trap_env_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "010UU"; -- 8..11: environment call from u/s/h/m
  -- RISC-V compliant asynchronous exceptions (interrupts) --
  constant trap_msi_c      : std_ulogic_vector(6 downto 0) := "1" & "0" & "00011"; -- 3:  machine software interrupt
  constant trap_mti_c      : std_ulogic_vector(6 downto 0) := "1" & "0" & "00111"; -- 7:  machine timer interrupt
  constant trap_mei_c      : std_ulogic_vector(6 downto 0) := "1" & "0" & "01011"; -- 11: machine external interrupt
  -- NEORV32-specific (RISC-V custom) asynchronous exceptions (interrupts) --
  constant trap_firq0_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10000"; -- 16: fast interrupt 0
  constant trap_firq1_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10001"; -- 17: fast interrupt 1
  constant trap_firq2_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10010"; -- 18: fast interrupt 2
  constant trap_firq3_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10011"; -- 19: fast interrupt 3
  constant trap_firq4_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10100"; -- 20: fast interrupt 4
  constant trap_firq5_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10101"; -- 21: fast interrupt 5
  constant trap_firq6_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10110"; -- 22: fast interrupt 6
  constant trap_firq7_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10111"; -- 23: fast interrupt 7
  constant trap_firq8_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "11000"; -- 24: fast interrupt 8
  constant trap_firq9_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "11001"; -- 25: fast interrupt 9
  constant trap_firq10_c   : std_ulogic_vector(6 downto 0) := "1" & "0" & "11010"; -- 26: fast interrupt 10
  constant trap_firq11_c   : std_ulogic_vector(6 downto 0) := "1" & "0" & "11011"; -- 27: fast interrupt 11
  constant trap_firq12_c   : std_ulogic_vector(6 downto 0) := "1" & "0" & "11100"; -- 28: fast interrupt 12
  constant trap_firq13_c   : std_ulogic_vector(6 downto 0) := "1" & "0" & "11101"; -- 29: fast interrupt 13
  constant trap_firq14_c   : std_ulogic_vector(6 downto 0) := "1" & "0" & "11110"; -- 30: fast interrupt 14
  constant trap_firq15_c   : std_ulogic_vector(6 downto 0) := "1" & "0" & "11111"; -- 31: fast interrupt 15
  -- entering debug mode (sync./async. exceptions) --
  constant trap_db_break_c : std_ulogic_vector(6 downto 0) := "0" & "1" & "00001"; -- 1: break instruction (sync)
  constant trap_db_trig_c  : std_ulogic_vector(6 downto 0) := "0" & "1" & "00010"; -- 2: hardware trigger (sync)
  constant trap_db_halt_c  : std_ulogic_vector(6 downto 0) := "1" & "1" & "00011"; -- 3: external halt request (async)
  constant trap_db_step_c  : std_ulogic_vector(6 downto 0) := "1" & "1" & "00100"; -- 4: single-stepping (async)

  -- Trap System ----------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- exception source bits --
  constant exc_iaccess_c  : natural :=  0; -- instruction access fault
  constant exc_illegal_c  : natural :=  1; -- illegal instruction
  constant exc_ialign_c   : natural :=  2; -- instruction address misaligned
  constant exc_ecall_c    : natural :=  3; -- environment call
  constant exc_ebreak_c   : natural :=  4; -- breakpoint
  constant exc_salign_c   : natural :=  5; -- store address misaligned
  constant exc_lalign_c   : natural :=  6; -- load address misaligned
  constant exc_saccess_c  : natural :=  7; -- store access fault
  constant exc_laccess_c  : natural :=  8; -- load access fault
  -- for debug mode only --
  constant exc_db_break_c : natural :=  9; -- enter debug mode via ebreak instruction
  constant exc_db_hw_c    : natural := 10; -- enter debug mode via hw trigger
  --
  constant exc_width_c    : natural := 11; -- length of this list in bits
  -- interrupt source bits --
  constant irq_msi_irq_c  : natural :=  0; -- machine software interrupt
  constant irq_mti_irq_c  : natural :=  1; -- machine timer interrupt
  constant irq_mei_irq_c  : natural :=  2; -- machine external interrupt
  constant irq_firq_0_c   : natural :=  3; -- fast interrupt channel 0
  constant irq_firq_1_c   : natural :=  4; -- fast interrupt channel 1
  constant irq_firq_2_c   : natural :=  5; -- fast interrupt channel 2
  constant irq_firq_3_c   : natural :=  6; -- fast interrupt channel 3
  constant irq_firq_4_c   : natural :=  7; -- fast interrupt channel 4
  constant irq_firq_5_c   : natural :=  8; -- fast interrupt channel 5
  constant irq_firq_6_c   : natural :=  9; -- fast interrupt channel 6
  constant irq_firq_7_c   : natural := 10; -- fast interrupt channel 7
  constant irq_firq_8_c   : natural := 11; -- fast interrupt channel 8
  constant irq_firq_9_c   : natural := 12; -- fast interrupt channel 9
  constant irq_firq_10_c  : natural := 13; -- fast interrupt channel 10
  constant irq_firq_11_c  : natural := 14; -- fast interrupt channel 11
  constant irq_firq_12_c  : natural := 15; -- fast interrupt channel 12
  constant irq_firq_13_c  : natural := 16; -- fast interrupt channel 13
  constant irq_firq_14_c  : natural := 17; -- fast interrupt channel 14
  constant irq_firq_15_c  : natural := 18; -- fast interrupt channel 15
  -- for debug mode only --
  constant irq_db_halt_c  : natural := 19; -- enter debug mode via external halt request
  constant irq_db_step_c  : natural := 20; -- enter debug mode via single-stepping
  --
  constant irq_width_c    : natural := 21; -- length of this list in bits

  -- Privilege Modes ------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant priv_mode_m_c : std_ulogic := '1'; -- machine mode
  constant priv_mode_u_c : std_ulogic := '0'; -- user mode

  -- HPM Event System -----------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant hpmcnt_event_cy_c          : natural := 0;  -- Active cycle
  constant hpmcnt_event_tm_c          : natural := 1;  -- Time (unused/reserved)
  constant hpmcnt_event_ir_c          : natural := 2;  -- Retired instruction
  --constant hpmcnt_event_cir_c       : natural := 3;  -- Retired compressed instruction
  --constant hpmcnt_event_wait_if_c   : natural := 4;  -- Instruction fetch memory wait cycle
  --constant hpmcnt_event_wait_ii_c   : natural := 5;  -- Instruction issue wait cycle
  --constant hpmcnt_event_wait_mc_c   : natural := 6;  -- Multi-cycle ALU-operation wait cycle
  --constant hpmcnt_event_load_c      : natural := 7;  -- Load operation
  --constant hpmcnt_event_store_c       : natural := 8;  -- Store operation
  --constant hpmcnt_event_wait_ls_c     : natural := 9;  -- Load/store memory wait cycle
  --constant hpmcnt_event_tbranch_c     : natural := 12; -- Conditional taken branch
  constant hpmcnt_event_ecc_se_imem   : natural := 3; -- Register file single error
  constant hpmcnt_event_ecc_de_imem   : natural := 4; -- Register file double error
  constant hpmcnt_event_ecc_se_dmem   : natural := 5; -- Data memory single error
  constant hpmcnt_event_ecc_de_dmem   : natural := 6; -- Data memory double error
  constant hpmcnt_event_ecc_se_regfile: natural := 7; -- Register file single error
  constant hpmcnt_event_ecc_de_regfile: natural := 8; -- Register file double error
  constant hpmcnt_event_iv            : natural := 9; -- Instruction validator detecting an error
  constant hpmcnt_event_jump_c        : natural := 10; -- Unconditional jump
  constant hpmcnt_event_branch_c      : natural := 11; -- Conditional branch (taken or not taken)
  constant hpmcnt_event_dsp_timeout   : natural := 12; -- One of the DSPs timed out
  constant hpmcnt_event_trap_c        : natural := 13; -- Entered trap
  constant hpmcnt_event_illegal_c     : natural := 14; -- Illegal instruction exception
  --
  constant hpmcnt_event_size_c    : natural := 15; -- length of this list

-- ****************************************************************************************************************************
-- Helper Functions
-- ****************************************************************************************************************************

  function index_size_f(input : natural) return natural;
  function cond_sel_int_f(cond : boolean; val_t : integer; val_f : integer) return integer;
  function cond_sel_natural_f(cond : boolean; val_t : natural; val_f : natural) return natural;
  function cond_sel_suv_f(cond : boolean; val_t : std_ulogic_vector; val_f : std_ulogic_vector) return std_ulogic_vector;
  function cond_sel_string_f(cond : boolean; val_t : string; val_f : string) return string;
  function bool_to_ulogic_f(cond : boolean) return std_ulogic;
  function bin_to_gray_f(input : std_ulogic_vector) return std_ulogic_vector;
  function gray_to_bin_f(input : std_ulogic_vector) return std_ulogic_vector;
  function or_reduce_f(input : std_ulogic_vector) return std_ulogic;
  function and_reduce_f(input : std_ulogic_vector) return std_ulogic;
  function xor_reduce_f(input : std_ulogic_vector) return std_ulogic;
  function su_undefined_f(input : std_ulogic) return boolean;
  function to_hexchar_f(input : std_ulogic_vector(3 downto 0)) return character;
  function to_hstring32_f(input : std_ulogic_vector(31 downto 0)) return string;
  function bit_rev_f(input : std_ulogic_vector) return std_ulogic_vector;
  function is_power_of_two_f(input : natural) return boolean;
  function bswap32_f(input : std_ulogic_vector) return std_ulogic_vector;
  function popcount_f(input : std_ulogic_vector) return natural;
  function leading_zeros_f(input : std_ulogic_vector) return natural;
  impure function mem32_init_f(init : mem32_t; depth : natural) return mem32_t;

-- ****************************************************************************************************************************
-- NEORV32 Processor Top Entity (component prototype)
-- ****************************************************************************************************************************

  component neorv32_top
    generic (
      -- General --
      CLOCK_FREQUENCY            : natural;
      HART_ID                    : std_ulogic_vector(31 downto 0) := x"00000000";
      VENDOR_ID                  : std_ulogic_vector(31 downto 0) := x"00000000";
      INT_BOOTLOADER_EN          : boolean := false;
      -- On-Chip Debugger (OCD) --
      ON_CHIP_DEBUGGER_EN        : boolean := false;
      DM_LEGACY_MODE             : boolean := false;
      -- RISC-V CPU Extensions --
      CPU_EXTENSION_RISCV_A      : boolean := false;
      CPU_EXTENSION_RISCV_B      : boolean := false;
      CPU_EXTENSION_RISCV_C      : boolean := false;
      CPU_EXTENSION_RISCV_E      : boolean := false;
      CPU_EXTENSION_RISCV_M      : boolean := false;
      CPU_EXTENSION_RISCV_U      : boolean := false;
      CPU_EXTENSION_RISCV_Zfinx  : boolean := false;
      CPU_EXTENSION_RISCV_Zicntr : boolean := true;
      CPU_EXTENSION_RISCV_Zihpm  : boolean := false;
      CPU_EXTENSION_RISCV_Zmmul  : boolean := false;
      CPU_EXTENSION_RISCV_Zxcfu  : boolean := false;
      -- Tuning Options --
      FAST_MUL_EN                : boolean := false;
      FAST_SHIFT_EN              : boolean := false;
      REGFILE_HW_RST             : boolean := false;
      -- Physical Memory Protection (PMP) --
      PMP_NUM_REGIONS            : natural range 0 to 16 := 0;
      PMP_MIN_GRANULARITY        : natural := 4;
      -- Hardware Performance Monitors (HPM) --
      HPM_NUM_CNTS               : natural range 0 to 13 := 0;
      HPM_CNT_WIDTH              : natural range 0 to 64 := 40;
      -- Atomic Memory Access - Reservation Set Granularity --
      AMO_RVS_GRANULARITY        : natural := 4;
      -- Internal Instruction memory (IMEM) --
      MEM_INT_IMEM_EN            : boolean := false;
      MEM_INT_IMEM_SIZE          : natural := 16*1024;
      MEM_INT_IMEM_PREFETCH      : boolean := false;
      MEM_INT_PREFETCH_BASE      : std_logic_vector(31 downto 0) := x"00000000";
      MEM_INT_IMEM_ECC_BP        : boolean := false;
      MEM_INT_IV_EN              : boolean := false;
      -- Internal Data memory (DMEM) --
      MEM_INT_DMEM_EN            : boolean := false;
      MEM_INT_DMEM_SIZE          : natural := 8*1024;
      -- Internal Instruction Cache (iCACHE) --
      ICACHE_EN                  : boolean                  := false;
      ICACHE_NUM_BLOCKS          : natural range 1 to 256   := 4;
      ICACHE_BLOCK_SIZE          : natural range 4 to 2**16 := 64;
      ICACHE_ASSOCIATIVITY       : natural range 1 to 2     := 1;
      -- Internal Data Cache (dCACHE) --
      DCACHE_EN                  : boolean                  := false;
      DCACHE_NUM_BLOCKS          : natural range 1 to 256   := 4;
      DCACHE_BLOCK_SIZE          : natural range 4 to 2**16 := 64;
      -- External memory interface (WISHBONE) --
      MEM_EXT_EN                 : boolean := false;
      MEM_EXT_TIMEOUT            : natural := 255;
      MEM_EXT_PIPE_MODE          : boolean := false;
      MEM_EXT_BIG_ENDIAN         : boolean := false;
      MEM_EXT_ASYNC_RX           : boolean := false;
      MEM_EXT_ASYNC_TX           : boolean := false;
      -- External Interrupts Controller (XIRQ) --
      XIRQ_NUM_CH                : natural range 0 to 32          := 0;
      XIRQ_TRIGGER_TYPE          : std_ulogic_vector(31 downto 0) := x"ffffffff";
      XIRQ_TRIGGER_POLARITY      : std_ulogic_vector(31 downto 0) := x"ffffffff";
      -- Processor peripherals --
      IO_GPIO_NUM                : natural range 0 to 64          := 0;
      IO_MTIME_EN                : boolean                        := false;
      IO_UART0_EN                : boolean                        := false;
      IO_UART0_RX_FIFO           : natural range 1 to 2**15       := 1;
      IO_UART0_TX_FIFO           : natural range 1 to 2**15       := 1;
      IO_UART1_EN                : boolean                        := false;
      IO_UART1_RX_FIFO           : natural range 1 to 2**15       := 1;
      IO_UART1_TX_FIFO           : natural range 1 to 2**15       := 1;
      IO_SPI_EN                  : boolean                        := false;
      IO_SPI_FIFO                : natural range 1 to 2**15       := 1;
      IO_SDI_EN                  : boolean                        := false;
      IO_SDI_FIFO                : natural range 1 to 2**15       := 1;
      IO_TWI_EN                  : boolean                        := false;
      IO_PWM_NUM_CH              : natural range 0 to 12          := 0;
      IO_WDT_EN                  : boolean                        := false;
      IO_TRNG_EN                 : boolean                        := false;
      IO_TRNG_FIFO               : natural range 1 to 2**15       := 1;
      IO_CFS_EN                  : boolean                        := false;
      IO_CFS_CONFIG              : std_ulogic_vector(31 downto 0) := x"00000000";
      IO_CFS_IN_SIZE             : natural                        := 32;
      IO_CFS_OUT_SIZE            : natural                        := 32;
      IO_NEOLED_EN               : boolean                        := false;
      IO_NEOLED_TX_FIFO          : natural range 1 to 2**15       := 1;
      IO_GPTMR_EN                : boolean                        := false;
      IO_XIP_EN                  : boolean                        := false;
      IO_ONEWIRE_EN              : boolean                        := false;
      IO_DMA_EN                  : boolean                        := false;
      IO_SLINK_EN                : boolean                        := false;
      IO_SLINK_RX_FIFO           : natural range 1 to 2**15       := 1;
      IO_SLINK_TX_FIFO           : natural range 1 to 2**15       := 1;
      IO_CRC_EN                  : boolean                        := false
    );
    port (
      -- Global control --
      clk_i          : in  std_ulogic;
      rstn_i         : in  std_ulogic;
      -- JTAG on-chip debugger interface --
      jtag_trst_i    : in  std_ulogic := 'U';
      jtag_tck_i     : in  std_ulogic := 'U';
      jtag_tdi_i     : in  std_ulogic := 'U';
      jtag_tdo_o     : out std_ulogic;
      jtag_tms_i     : in  std_ulogic := 'U';
      -- Wishbone bus interface (available if MEM_EXT_EN = true) --
      wb_tag_o       : out std_ulogic_vector(02 downto 0);
      wb_adr_o       : out std_ulogic_vector(31 downto 0);
      wb_dat_i       : in  std_ulogic_vector(31 downto 0) := (others => 'U');
      wb_dat_o       : out std_ulogic_vector(31 downto 0);
      wb_we_o        : out std_ulogic;
      wb_sel_o       : out std_ulogic_vector(03 downto 0);
      wb_stb_o       : out std_ulogic;
      wb_cyc_o       : out std_ulogic;
      wb_ack_i       : in  std_ulogic := 'L';
      wb_err_i       : in  std_ulogic := 'L';
      -- Stream Link Interface (available if IO_SLINK_EN = true) --
      slink_rx_dat_i : in  std_ulogic_vector(31 downto 0) := (others => 'U');
      slink_rx_val_i : in  std_ulogic := 'L';
      slink_rx_rdy_o : out std_ulogic;
      slink_tx_dat_o : out std_ulogic_vector(31 downto 0);
      slink_tx_val_o : out std_ulogic;
      slink_tx_rdy_i : in  std_ulogic := 'L';
      -- Advanced memory control signals --
      fence_o        : out std_ulogic;
      fencei_o       : out std_ulogic;
      -- XIP (execute in place via SPI) signals (available if IO_XIP_EN = true) --
      xip_csn_o      : out std_ulogic;
      xip_clk_o      : out std_ulogic;
      xip_dat_i      : in  std_ulogic := 'L';
      xip_dat_o      : out std_ulogic;
      -- GPIO (available if IO_GPIO_NUM > 0) --
      gpio_o         : out std_ulogic_vector(63 downto 0);
      gpio_i         : in  std_ulogic_vector(63 downto 0) := (others => 'U');
      -- primary UART0 (available if IO_UART0_EN = true) --
      uart0_txd_o    : out std_ulogic;
      uart0_rxd_i    : in  std_ulogic := 'U';
      uart0_rts_o    : out std_ulogic;
      uart0_cts_i    : in  std_ulogic := 'L';
      -- secondary UART1 (available if IO_UART1_EN = true) --
      uart1_txd_o    : out std_ulogic;
      uart1_rxd_i    : in  std_ulogic := 'U'; -- UART1 receive data
      uart1_rts_o    : out std_ulogic;
      uart1_cts_i    : in  std_ulogic := 'L';
      -- SPI (available if IO_SPI_EN = true) --
      spi_clk_o      : out std_ulogic;
      spi_dat_o      : out std_ulogic;
      spi_dat_i      : in  std_ulogic := 'U';
      spi_csn_o      : out std_ulogic_vector(07 downto 0); -- SPI CS
      -- SDI (available if IO_SDI_EN = true) --
      sdi_clk_i      : in  std_ulogic := 'U';
      sdi_dat_o      : out std_ulogic;
      sdi_dat_i      : in  std_ulogic := 'U';
      sdi_csn_i      : in  std_ulogic := 'H';
      -- TWI (available if IO_TWI_EN = true) --
      twi_sda_i      : in  std_ulogic := 'H';
      twi_sda_o      : out std_ulogic;
      twi_scl_i      : in  std_ulogic := 'H';
      twi_scl_o      : out std_ulogic;
      -- 1-Wire Interface (available if IO_ONEWIRE_EN = true) --
      onewire_i      : in  std_ulogic := 'H';
      onewire_o      : out std_ulogic;
      -- PWM (available if IO_PWM_NUM_CH > 0) --
      pwm_o          : out std_ulogic_vector(11 downto 0); -- pwm channels
      -- Custom Functions Subsystem IO --
      cfs_in_i       : in  std_ulogic_vector(IO_CFS_IN_SIZE-1 downto 0) := (others => 'U');
      cfs_out_o      : out std_ulogic_vector(IO_CFS_OUT_SIZE-1 downto 0);
      -- NeoPixel-compatible smart LED interface (available if IO_NEOLED_EN = true) --
      neoled_o       : out std_ulogic;
      -- External platform interrupts (available if XIRQ_NUM_CH > 0) --
      xirq_i         : in  std_ulogic_vector(31 downto 0) := (others => 'L');
      -- CPU Interrupts --
      mtime_irq_i    : in  std_ulogic := 'L';
      msw_irq_i      : in  std_ulogic := 'L';
      mext_irq_i     : in  std_ulogic := 'L'
    );
  end component;

end neorv32_package;

package body neorv32_package is

-- ****************************************************************************************************************************
-- Functions
-- ****************************************************************************************************************************

  -- Minimal required number of bits to represent <input> numbers ---------------------------
  -- -------------------------------------------------------------------------------------------
  function index_size_f(input : natural) return natural is
  begin
    for i in 0 to natural'high loop
      if (2**i >= input) then
        return i;
      end if;
    end loop;
    return 0;
  end function index_size_f;

  -- Conditional select integer -------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function cond_sel_int_f(cond : boolean; val_t : integer; val_f : integer) return integer is
  begin
    if (cond = true) then
      return val_t;
    else
      return val_f;
    end if;
  end function cond_sel_int_f;

  -- Conditional select natural -------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function cond_sel_natural_f(cond : boolean; val_t : natural; val_f : natural) return natural is
  begin
    if (cond = true) then
      return val_t;
    else
      return val_f;
    end if;
  end function cond_sel_natural_f;

  -- Conditional select std_ulogic_vector ---------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function cond_sel_suv_f(cond : boolean; val_t : std_ulogic_vector; val_f : std_ulogic_vector) return std_ulogic_vector is
  begin
    if (cond = true) then
      return val_t;
    else
      return val_f;
    end if;
  end function cond_sel_suv_f;

  -- Conditional select string --------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function cond_sel_string_f(cond : boolean; val_t : string; val_f : string) return string is
  begin
    if (cond = true) then
      return val_t;
    else
      return val_f;
    end if;
  end function cond_sel_string_f;

  -- Convert boolean to std_ulogic ----------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function bool_to_ulogic_f(cond : boolean) return std_ulogic is
  begin
    if (cond = true) then
      return '1';
    else
      return '0';
    end if;
  end function bool_to_ulogic_f;

  -- Convert binary to gray -----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function bin_to_gray_f(input : std_ulogic_vector) return std_ulogic_vector is
    variable tmp_v : std_ulogic_vector(input'range);
  begin
    tmp_v(input'length-1) := input(input'length-1); -- keep MSB
    for i in input'length-2 downto 0 loop
      tmp_v(i) := input(i) xor input(i+1);
    end loop;
    return tmp_v;
  end function bin_to_gray_f;

  -- Convert gray to binary -----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function gray_to_bin_f(input : std_ulogic_vector) return std_ulogic_vector is
    variable tmp_v : std_ulogic_vector(input'range);
  begin
    tmp_v(input'length-1) := input(input'length-1); -- keep MSB
    for i in input'length-2 downto 0 loop
      tmp_v(i) := tmp_v(i+1) xor input(i);
    end loop;
    return tmp_v;
  end function gray_to_bin_f;

  -- OR all bits ----------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function or_reduce_f(input : std_ulogic_vector) return std_ulogic is
    variable tmp_v : std_ulogic;
  begin
    tmp_v := '0';
    for i in input'range loop
      tmp_v := tmp_v or input(i);
    end loop;
    return tmp_v;
  end function or_reduce_f;

  -- AND all bits ---------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function and_reduce_f(input : std_ulogic_vector) return std_ulogic is
    variable tmp_v : std_ulogic;
  begin
    tmp_v := '1';
    for i in input'range loop
      tmp_v := tmp_v and input(i);
    end loop;
    return tmp_v;
  end function and_reduce_f;

  -- XOR all bits ---------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function xor_reduce_f(input : std_ulogic_vector) return std_ulogic is
    variable tmp_v : std_ulogic;
  begin
    tmp_v := '0';
    for i in input'range loop
      tmp_v := tmp_v xor input(i);
    end loop;
    return tmp_v;
  end function xor_reduce_f;

  -- Check if std_ulogic is not '1' or '0' --------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function su_undefined_f(input : std_ulogic) return boolean is
  begin
    case input is
      when '1' | '0' => return false;
      when others    => return true;
    end case;
  end function su_undefined_f;

  -- Convert std_ulogic_vector to lowercase HEX char ----------------------------------------
  -- -------------------------------------------------------------------------------------------
  function to_hexchar_f(input : std_ulogic_vector(3 downto 0)) return character is
    variable hex_v : string(1 to 16);
  begin
    hex_v := "0123456789abcdef";
    if (su_undefined_f(input(3)) = true) or (su_undefined_f(input(2)) = true) or
       (su_undefined_f(input(1)) = true) or (su_undefined_f(input(0)) = true) then
      return '?';
    else
      return hex_v(to_integer(unsigned(input)) + 1);
    end if;
  end function to_hexchar_f;

  -- Convert 32-bit std_ulogic_vector to hex string -----------------------------------------
  -- -------------------------------------------------------------------------------------------
  function to_hstring32_f(input : std_ulogic_vector(31 downto 0)) return string is
    variable res_v : string(1 to 8);
  begin
    for i in 7 downto 0 loop
      res_v(8-i) := to_hexchar_f(input(i*4+3 downto i*4+0));
    end loop;
    return res_v;
  end function to_hstring32_f;

  -- Bit reversal ---------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function bit_rev_f(input : std_ulogic_vector) return std_ulogic_vector is
    variable output_v : std_ulogic_vector(input'range);
  begin
    for i in 0 to input'length-1 loop
      output_v(input'length-i-1) := input(i);
    end loop;
    return output_v;
  end function bit_rev_f;

  -- Test if input number is a power of two -------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function is_power_of_two_f(input : natural) return boolean is
    variable tmp : unsigned(31 downto 0);
  begin
    if (input = 0) then
      return false;
    elsif (input = 1) then
      return true;
    else
      tmp := to_unsigned(input, 32);
      if ((tmp and (tmp - 1)) = 0) then
        return true;
      else
        return false;
      end if;
    end if;
  end function is_power_of_two_f;

  -- Swap all bytes of a 32-bit word (endianness conversion) --------------------------------
  -- -------------------------------------------------------------------------------------------
  function bswap32_f(input : std_ulogic_vector) return std_ulogic_vector is
    variable output_v : std_ulogic_vector(input'range);
  begin
    output_v(07 downto 00) := input(31 downto 24);
    output_v(15 downto 08) := input(23 downto 16);
    output_v(23 downto 16) := input(15 downto 08);
    output_v(31 downto 24) := input(07 downto 00);
    return output_v;
  end function bswap32_f;

  -- Population count (number of set bits) --------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function popcount_f(input : std_ulogic_vector) return natural is
    variable cnt_v : natural range 0 to input'length;
  begin
    cnt_v := 0;
    for i in input'length-1 downto 0 loop
      if (input(i) = '1') then
        cnt_v := cnt_v + 1;
      end if;
    end loop;
    return cnt_v;
  end function popcount_f;

  -- Count leading zeros --------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function leading_zeros_f(input : std_ulogic_vector) return natural is
    variable cnt_v : natural range 0 to input'length;
  begin
    cnt_v := 0;
    for i in input'length-1 downto 0 loop
      if (input(i) = '0') then
        cnt_v := cnt_v + 1;
      else
        exit;
      end if;
    end loop;
    return cnt_v;
  end function leading_zeros_f;

  -- Initialize mem32_t array from another mem32_t array ------------------------------------
  -- -------------------------------------------------------------------------------------------
  impure function mem32_init_f(init : mem32_t; depth : natural) return mem32_t is
    variable mem_v : mem32_t(0 to depth-1);
  begin
    mem_v := (others => (others => '0')); -- [IMPORTANT] make sure remaining memory entries are set to zero
    if (init'length > depth) then
      return mem_v;
    end if;
    for i in 0 to init'length-1 loop -- initialize only in range of source data array
      mem_v(i) := init(i);
    end loop;
    return mem_v;
  end function mem32_init_f;


end neorv32_package;

-- ****************************************************************************************************************************
-- Additional Packages
-- ****************************************************************************************************************************

  -- Prototype Definition: bootloader_init_image --------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- > memory content in 'neorv32_bootloader_image.vhd', auto-generated by 'image_gen'
  -- > used by 'neorv32_boot_rom.vhd'
  -- > enables body-only recompile in case of firmware change (NEORV32 PR #338)

library ieee;
use ieee.std_logic_1164.all;

library neorv32;
use neorv32.neorv32_package.all;

package neorv32_bootloader_image is
  constant bootloader_init_image : mem32_t;
end neorv32_bootloader_image;


  -- Prototype Definition: neorv32_application_image ----------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- > memory content in 'neorv32_application_image.vhd', auto-generated by 'image_gen'
  -- > used by 'mem/neorv32_imem.*.vhd'
  -- > enables body-only recompile in case of firmware change (NEORV32 PR #338)

library ieee;
use ieee.std_logic_1164.all;

library neorv32;
use neorv32.neorv32_package.all;

package neorv32_application_image is
  constant application_init_image : mem32_t := (
x"de067139",
x"0080dc22",
x"fca42623",
x"152387ae",
x"1723fcf4",
x"1623fe04",
x"1523fe04",
x"2783fe04",
x"53dcfcc4",
x"fef42223",
x"fcc42783",
x"0047d783",
x"fcf41e23",
x"fca45783",
x"fcf41923",
x"fc041f23",
x"5783a221",
x"f793fde4",
x"07c20ff7",
x"182387c1",
x"0793fcf4",
x"85befd04",
x"fe442503",
x"2a232ad5",
x"2503fca4",
x"24b5fe44",
x"fea42223",
x"fd442783",
x"5783eb95",
x"0785fea4",
x"fef41523",
x"fe442783",
x"43dc439c",
x"00079783",
x"07c287a1",
x"07c287c1",
x"8b8583c1",
x"83c107c2",
x"fee45703",
x"172397ba",
x"a89dfef4",
x"fec45783",
x"16230785",
x"2783fef4",
x"43dcfd44",
x"00079783",
x"83c107c2",
x"c39d8b85",
x"fd442783",
x"978343dc",
x"87a50007",
x"87c107c2",
x"83c107c2",
x"07c28b85",
x"570383c1",
x"97bafee4",
x"fef41723",
x"fd442783",
x"c79d439c",
x"fd442783",
x"2023439c",
x"2783fef4",
x"4398fe04",
x"fd442783",
x"2783c398",
x"4398fe44",
x"fe042783",
x"2783c398",
x"2703fe44",
x"c398fe04",
x"fd241783",
x"0007cd63",
x"fd241783",
x"83c107c2",
x"07c20785",
x"07c283c1",
x"192387c1",
x"1783fcf4",
x"07c2fde4",
x"078583c1",
x"83c107c2",
x"fcf41f23",
x"fde41703",
x"fdc41783",
x"eef749e3",
x"fec45783",
x"07c2078a",
x"570383c1",
x"8f99fea4",
x"83c107c2",
x"fee45703",
x"172397ba",
x"1783fef4",
x"5b63fca4",
x"260300f0",
x"0593fcc4",
x"25035660",
x"2c25fe44",
x"fea42223",
x"fe442783",
x"853e439c",
x"2c232251",
x"0793fca4",
x"85befd04",
x"fe442503",
x"20232075",
x"2783fea4",
x"eb95fe04",
x"fe442783",
x"2023439c",
x"a025fef4",
x"fe442783",
x"978343dc",
x"57030007",
x"85bafee4",
x"00ef853e",
x"87aa4050",
x"fef41723",
x"fe042783",
x"2023439c",
x"2783fef4",
x"fbf9fe04",
x"fe442783",
x"85be439c",
x"fd842503",
x"2c232aad",
x"4601fca4",
x"5b400593",
x"fe442503",
x"22232a6d",
x"2783fea4",
x"439cfe44",
x"fef42023",
x"2783a025",
x"43dcfe44",
x"00079783",
x"fee45703",
x"853e85ba",
x"3ab000ef",
x"172387aa",
x"2783fef4",
x"439cfe04",
x"fef42023",
x"fe042783",
x"5783fbf9",
x"853efee4",
x"546250f2",
x"80826121",
x"ce221101",
x"26231000",
x"2423fea4",
x"2783feb4",
x"9783fe84",
x"ce630027",
x"a0310207",
x"fec42783",
x"2623439c",
x"2783fef4",
x"cf81fec4",
x"fec42783",
x"970343dc",
x"27830027",
x"9783fe84",
x"1fe30027",
x"2783fcf7",
x"a815fec4",
x"fec42783",
x"2623439c",
x"2783fef4",
x"c385fec4",
x"fec42783",
x"978343dc",
x"07c20007",
x"f79383c1",
x"27030ff7",
x"1703fe84",
x"9be30007",
x"2783fce7",
x"853efec4",
x"61054472",
x"71798082",
x"1800d622",
x"fca42e23",
x"fe042623",
x"2783a01d",
x"439cfdc4",
x"fef42423",
x"fdc42783",
x"fec42703",
x"2783c398",
x"2623fdc4",
x"2783fef4",
x"2e23fe84",
x"2783fcf4",
x"ffe1fdc4",
x"fec42783",
x"5432853e",
x"80826145",
x"d6227179",
x"2e231800",
x"2783fca4",
x"439cfdc4",
x"fef42623",
x"fdc42783",
x"242343dc",
x"2783fef4",
x"43d8fec4",
x"fdc42783",
x"2783c3d8",
x"2703fec4",
x"c3d8fe84",
x"fdc42783",
x"4398439c",
x"fdc42783",
x"2783c398",
x"a023fec4",
x"27830007",
x"853efec4",
x"61455432",
x"71798082",
x"1800d622",
x"fca42e23",
x"fcb42c23",
x"fdc42783",
x"262343dc",
x"2783fef4",
x"43d8fd84",
x"fdc42783",
x"2783c3d8",
x"2703fd84",
x"c3d8fec4",
x"fd842783",
x"27834398",
x"c398fdc4",
x"fd842783",
x"fdc42703",
x"2783c398",
x"853efdc4",
x"61455432",
x"715d8082",
x"c4a2c686",
x"2e230880",
x"2c23faa4",
x"2a23fab4",
x"4785fac4",
x"fcf42e23",
x"fbc42783",
x"fef42623",
x"fa042e23",
x"fe042023",
x"fc042c23",
x"2783a291",
x"0785fd84",
x"fcf42c23",
x"fec42783",
x"fef42423",
x"fc042a23",
x"fc042623",
x"2783a01d",
x"0785fd44",
x"fcf42a23",
x"fe842783",
x"2423439c",
x"2783fef4",
x"cf89fe84",
x"fcc42783",
x"26230785",
x"2703fcf4",
x"2783fcc4",
x"4ae3fdc4",
x"a011fcf7",
x"27830001",
x"2823fdc4",
x"a0f1fcf4",
x"fd442783",
x"2783e385",
x"2223fe84",
x"2783fef4",
x"439cfe84",
x"fef42423",
x"fd042783",
x"282317fd",
x"a059fcf4",
x"fd042783",
x"2783c781",
x"e385fe84",
x"fec42783",
x"fef42223",
x"fec42783",
x"2623439c",
x"2783fef4",
x"17fdfd44",
x"fcf42a23",
x"2783a8b1",
x"43d8fec4",
x"fe842783",
x"278343d4",
x"2603fb84",
x"85b6fb44",
x"9782853a",
x"416387aa",
x"278302f0",
x"2223fec4",
x"2783fef4",
x"439cfec4",
x"fef42623",
x"fd442783",
x"2a2317fd",
x"a839fcf4",
x"fe842783",
x"fef42223",
x"fe842783",
x"2423439c",
x"2783fef4",
x"17fdfd04",
x"fcf42823",
x"fe042783",
x"2783c799",
x"2703fe04",
x"c398fe44",
x"2783a029",
x"2e23fe44",
x"2783faf4",
x"2023fe44",
x"2783fef4",
x"49e3fd44",
x"2783f2f0",
x"5563fd04",
x"278300f0",
x"f38dfe84",
x"fe842783",
x"fef42623",
x"fec42783",
x"ea079de3",
x"fe042783",
x"0007a023",
x"fd842703",
x"c5634785",
x"278300e7",
x"a039fbc4",
x"fdc42783",
x"2e230786",
x"bdbdfcf4",
x"40b6853e",
x"61614426",
x"71798082",
x"d422d606",
x"2e231800",
x"2c23fca4",
x"2a23fcb4",
x"2783fcc4",
x"2583fdc4",
x"853efd44",
x"87aa28d9",
x"fef41723",
x"fd842783",
x"fd442583",
x"20d1853e",
x"162387aa",
x"1703fef4",
x"1783fee4",
x"07b3fec4",
x"853e40f7",
x"542250b2",
x"80826145",
x"ce221101",
x"26231000",
x"2423fea4",
x"2223feb4",
x"2783fec4",
x"ebadfe44",
x"fec42783",
x"00079783",
x"f007f793",
x"01079713",
x"27838741",
x"9783fec4",
x"07c20007",
x"83a183c1",
x"83c107c2",
x"87c107c2",
x"97138fd9",
x"87410107",
x"fec42783",
x"00e79023",
x"fe842783",
x"00079783",
x"f007f793",
x"01079713",
x"27838741",
x"9783fe84",
x"07c20007",
x"83a183c1",
x"83c107c2",
x"87c107c2",
x"97138fd9",
x"87410107",
x"fe842783",
x"00e79023",
x"fec42783",
x"00279783",
x"2783873e",
x"9783fe84",
x"07b30027",
x"853e40f7",
x"61054472",
x"71798082",
x"d422d606",
x"2e231800",
x"2c23fca4",
x"2783fcb4",
x"d783fdc4",
x"15230007",
x"1783fef4",
x"879dfea4",
x"87c107c2",
x"0ff7f793",
x"04a38b85",
x"4783fef4",
x"cb81fe94",
x"fea45783",
x"07f7f793",
x"87c107c2",
x"5783aa2d",
x"8b9dfea4",
x"fef41323",
x"fea41783",
x"07c2878d",
x"8bbd87c1",
x"fef41623",
x"fec45783",
x"07c20792",
x"570387c1",
x"8fd9fec4",
x"fef41623",
x"fe641783",
x"4705c789",
x"06e78163",
x"1703a861",
x"0793fec4",
x"c6630210",
x"079300e7",
x"16230220",
x"2783fef4",
x"4f88fd84",
x"fd842783",
x"27834bcc",
x"9603fd84",
x"27830007",
x"9683fd84",
x"27830027",
x"d783fd84",
x"17030387",
x"26c5fec4",
x"172387aa",
x"2783fef4",
x"d783fd84",
x"ebb103e7",
x"fee45703",
x"fd842783",
x"02e79f23",
x"2783a099",
x"8713fd84",
x"27830287",
x"d683fd84",
x"17830387",
x"8636fec4",
x"853a85be",
x"87aa2605",
x"fef41723",
x"fd842783",
x"03c7d783",
x"5703ef99",
x"2783fee4",
x"9e23fd84",
x"a80102e7",
x"fea45783",
x"fef41723",
x"0001a021",
x"0001a011",
x"fee45703",
x"fd842783",
x"0387d783",
x"853a85be",
x"87aa2d8d",
x"2783873e",
x"9c23fd84",
x"578302e7",
x"f793fee4",
x"172307f7",
x"5783fef4",
x"f793fea4",
x"07c2f007",
x"e79387c1",
x"07c20807",
x"570387c1",
x"8fd9fee4",
x"01079713",
x"27838741",
x"9023fdc4",
x"178300e7",
x"853efee4",
x"542250b2",
x"80826145",
x"d6067179",
x"1800d422",
x"fca42e23",
x"fdc42783",
x"fef42423",
x"fe842783",
x"22234fdc",
x"2783fef4",
x"9c23fe84",
x"27830207",
x"9d23fe84",
x"27830207",
x"9e23fe84",
x"27830207",
x"9f23fe84",
x"26230207",
x"a8bdfe04",
x"25034585",
x"f0effe84",
x"87aafd6f",
x"fef41123",
x"fe842783",
x"0387d703",
x"fe245783",
x"853e85ba",
x"87aa2b7d",
x"2783873e",
x"9c23fe84",
x"55fd02e7",
x"fe842503",
x"fa8ff0ef",
x"112387aa",
x"2783fef4",
x"d703fe84",
x"57830387",
x"85bafe24",
x"2b41853e",
x"873e87aa",
x"fe842783",
x"02e79c23",
x"fec42783",
x"2783eb89",
x"d703fe84",
x"27830387",
x"9d23fe84",
x"278302e7",
x"0785fec4",
x"fef42623",
x"fec42703",
x"fe442783",
x"f6f76ee3",
x"853e4781",
x"542250b2",
x"80826145",
x"de227139",
x"26230080",
x"2423fca4",
x"2223fcb4",
x"2023fcc4",
x"2023fcd4",
x"4785fe04",
x"fef42623",
x"fe042423",
x"fe042223",
x"fc442783",
x"4785e38d",
x"fcf42223",
x"2783a829",
x"0785fe84",
x"fef42423",
x"fe842783",
x"02f787b3",
x"2223078e",
x"2703fef4",
x"2783fe44",
x"60e3fcc4",
x"2783fef7",
x"17fdfe84",
x"fef42023",
x"fc842783",
x"9bf117fd",
x"2e230791",
x"2783fcf4",
x"87b3fe04",
x"078602f7",
x"fdc42703",
x"2c2397ba",
x"2423fcf4",
x"a8e9fe04",
x"fe042223",
x"2703a87d",
x"2783fec4",
x"0733fc44",
x"579302f7",
x"83c141f7",
x"00f706b3",
x"177d6741",
x"07b38f75",
x"222340f7",
x"2783fcf4",
x"9713fc44",
x"83410107",
x"fec42783",
x"83c107c2",
x"07c297ba",
x"1b2383c1",
x"2703fcf4",
x"2783fe84",
x"0733fe04",
x"278302f7",
x"97bafe44",
x"27030786",
x"97bafd84",
x"fd645703",
x"00e79023",
x"fec42783",
x"01079713",
x"57838341",
x"97bafd64",
x"83c107c2",
x"fcf41b23",
x"fd645783",
x"0ff7f793",
x"fcf41b23",
x"fe842703",
x"fe042783",
x"02f70733",
x"fe442783",
x"078697ba",
x"fdc42703",
x"570397ba",
x"9023fd64",
x"278300e7",
x"0785fec4",
x"fef42623",
x"fe442783",
x"22230785",
x"2703fef4",
x"2783fe44",
x"6ee3fe04",
x"2783f2f7",
x"0785fe84",
x"fef42423",
x"fe842703",
x"fe042783",
x"f2f760e3",
x"fc042783",
x"fdc42703",
x"2783c3d8",
x"2703fc04",
x"c798fd84",
x"fe042783",
x"02f787b3",
x"27030786",
x"97bafd84",
x"9bf117fd",
x"873e0791",
x"fc042783",
x"2703c7d8",
x"2783fe04",
x"c398fc04",
x"fe042783",
x"5472853e",
x"80826121",
x"de067139",
x"0080dc22",
x"fca42623",
x"873287ae",
x"fcf41523",
x"142387ba",
x"2783fcf4",
x"439cfcc4",
x"fef42623",
x"fcc42783",
x"242347dc",
x"2783fef4",
x"43dcfcc4",
x"fef42223",
x"fcc42783",
x"2023479c",
x"5783fef4",
x"1f23fca4",
x"1783fcf4",
x"873efde4",
x"fe042683",
x"fe442603",
x"fe842583",
x"fec42503",
x"3e4090ef",
x"873e87aa",
x"fc845783",
x"853a85be",
x"87aa2ccd",
x"fcf41423",
x"fc845783",
x"50f2853e",
x"61215462",
x"71598082",
x"d4a2d686",
x"2e231880",
x"2c23f8a4",
x"85b2f8b4",
x"86ba8636",
x"87ae873e",
x"f8f41b23",
x"1a2387b2",
x"87b6f8f4",
x"f8f41923",
x"182387ba",
x"2783f8f4",
x"2023f984",
x"2623faf4",
x"a81dfe04",
x"fec42783",
x"17c1078a",
x"aa2397a2",
x"2783fa07",
x"078afec4",
x"97a217c1",
x"fb47a703",
x"fec42783",
x"17c1078a",
x"aa2397a2",
x"2783fce7",
x"0785fec4",
x"fef42623",
x"fec42703",
x"f3e3479d",
x"a81dfce7",
x"fa440713",
x"fa040793",
x"853e85ba",
x"2f00a0ef",
x"fea42223",
x"fe442783",
x"17c1078a",
x"a78397a2",
x"8713fd47",
x"27830017",
x"078afe44",
x"97a217c1",
x"fce7aa23",
x"fa042783",
x"0007c783",
x"2783f3f1",
x"2023f984",
x"a83dfaf4",
x"fa042783",
x"0007c703",
x"02c00793",
x"02f70163",
x"fa042783",
x"0007c683",
x"f9645783",
x"0ff7f713",
x"fa042783",
x"77138f35",
x"80230ff7",
x"270300e7",
x"1783fa04",
x"97baf924",
x"faf42023",
x"f9842703",
x"f9c42783",
x"2783973e",
x"ebe3fa04",
x"2783fae7",
x"2023f984",
x"a81dfaf4",
x"fa440713",
x"fa040793",
x"853e85ba",
x"2500a0ef",
x"fea42423",
x"fe842783",
x"17c1078a",
x"a78397a2",
x"8713fd47",
x"27830017",
x"078afe84",
x"97a217c1",
x"fce7aa23",
x"fa042783",
x"0007c783",
x"2783f3f1",
x"2023f984",
x"a83dfaf4",
x"fa042783",
x"0007c703",
x"02c00793",
x"02f70163",
x"fa042783",
x"0007c683",
x"f9445783",
x"0ff7f713",
x"fa042783",
x"77138f35",
x"80230ff7",
x"270300e7",
x"1783fa04",
x"97baf924",
x"faf42023",
x"f9842703",
x"f9c42783",
x"2783973e",
x"ebe3fa04",
x"2623fae7",
x"a0a1fe04",
x"fec42783",
x"17c1078a",
x"a78397a2",
x"5703fd47",
x"85baf904",
x"2a59853e",
x"182387aa",
x"2783f8f4",
x"078afec4",
x"97a217c1",
x"fb47a783",
x"f9045703",
x"853e85ba",
x"87aa2aa5",
x"f8f41823",
x"fec42783",
x"26230785",
x"2703fef4",
x"479dfec4",
x"fae7fae3",
x"f9045783",
x"50b6853e",
x"61655426",
x"71798082",
x"1800d622",
x"872e87aa",
x"fcf40fa3",
x"1e2387ba",
x"07a3fcf4",
x"06a3fe04",
x"0723fe04",
x"07a3fe04",
x"a069fe04",
x"fdc45783",
x"01879713",
x"07838761",
x"8fb9fdf4",
x"87e107e2",
x"0ff7f793",
x"06a38b85",
x"4783fef4",
x"8385fdf4",
x"fcf40fa3",
x"fed44703",
x"1e634785",
x"578300f7",
x"873efdc4",
x"07896791",
x"1e238fb9",
x"4785fcf4",
x"fef40723",
x"0723a019",
x"5783fe04",
x"8385fdc4",
x"fcf41e23",
x"fee44783",
x"5783cb89",
x"873efdc4",
x"8fd977e1",
x"fcf41e23",
x"5783a809",
x"873efdc4",
x"17fd67a1",
x"1e238ff9",
x"4783fcf4",
x"0785fef4",
x"fef407a3",
x"fef44703",
x"f9e3479d",
x"5783f6e7",
x"853efdc4",
x"61455432",
x"11018082",
x"cc22ce06",
x"87aa1000",
x"1723872e",
x"87bafef4",
x"fef41623",
x"fee45783",
x"fec45703",
x"853e85ba",
x"87aa2039",
x"40f2853e",
x"61054462",
x"11018082",
x"cc22ce06",
x"87aa1000",
x"1723872e",
x"87bafef4",
x"fef41623",
x"fee45783",
x"0ff7f793",
x"fec45703",
x"853e85ba",
x"87aa35dd",
x"fef41623",
x"fee45783",
x"07c283a1",
x"f79383c1",
x"57030ff7",
x"85bafec4",
x"35e1853e",
x"162387aa",
x"5783fef4",
x"853efec4",
x"446240f2",
x"80826105",
x"ce061101",
x"1000cc22",
x"fea42623",
x"152387ae",
x"2783fef4",
x"07c2fec4",
x"570387c1",
x"85bafea4",
x"3f91853e",
x"152387aa",
x"2783fef4",
x"83c1fec4",
x"87c107c2",
x"fea45703",
x"853e85ba",
x"87aa3f2d",
x"fef41523",
x"fea45783",
x"40f2853e",
x"61054462",
x"00008082",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"7fff9197",
x"86818193",
x"00000013",
x"00000013",
x"58818113",
x"ff017113",
x"00000297",
x"14c28293",
x"30529073",
x"00000097",
x"0d208093",
x"00008563",
x"00ef9082",
x"25730240",
x"4581f140",
x"30ef4601",
x"02971ba0",
x"82930000",
x"907300c2",
x"23033052",
x"bff50000",
x"32970000",
x"82930000",
x"83173f22",
x"03137fff",
x"8397fa23",
x"83937fff",
x"8c6300e3",
x"5a630062",
x"a5030073",
x"02910002",
x"00a32023",
x"4ae30311",
x"8082fe73",
x"b37346a1",
x"76133006",
x"ee110035",
x"99f1058d",
x"ca634e11",
x"238301c5",
x"20230005",
x"05110075",
x"48e315f1",
x"1073feb0",
x"80823003",
x"b37346a1",
x"42913006",
x"0055c563",
x"00357613",
x"0023ca11",
x"05050005",
x"47e315fd",
x"1073feb0",
x"80823003",
x"00052023",
x"15f10511",
x"fcb04ee3",
x"30031073",
x"20238082",
x"03110003",
x"fe734de3",
x"84068082",
x"ffff8297",
x"f0928293",
x"04028163",
x"ffff8297",
x"efc28293",
x"f14027f3",
x"b07346a1",
x"830a3006",
x"ffff8397",
x"2e838393",
x"0363938a",
x"37d10073",
x"00579d63",
x"7fff8317",
x"ed430313",
x"7fff8397",
x"f4038393",
x"00730363",
x"8317376d",
x"03137fff",
x"9397f363",
x"83937fff",
x"57638a43",
x"20230073",
x"03110003",
x"fe734de3",
x"808280a2",
x"342022f3",
x"34102373",
x"343023f3",
x"0000bfd5",
x"10210000",
x"30632042",
x"50a54084",
x"70e760c6",
x"91298108",
x"b16ba14a",
x"d1adc18c",
x"f1efe1ce",
x"02101231",
x"22523273",
x"429452b5",
x"62d672f7",
x"83189339",
x"a35ab37b",
x"c39cd3bd",
x"e3def3ff",
x"34432462",
x"14010420",
x"74c764e6",
x"548544a4",
x"b54ba56a",
x"95098528",
x"f5cfe5ee",
x"d58dc5ac",
x"26723653",
x"06301611",
x"66f676d7",
x"46b45695",
x"a77ab75b",
x"87389719",
x"e7fef7df",
x"c7bcd79d",
x"58e548c4",
x"78a76886",
x"18610840",
x"38232802",
x"d9edc9cc",
x"f9afe98e",
x"99698948",
x"b92ba90a",
x"4ad45af5",
x"6a967ab7",
x"0a501a71",
x"2a123a33",
x"cbdcdbfd",
x"eb9efbbf",
x"8b589b79",
x"ab1abb3b",
x"7c876ca6",
x"5cc54ce4",
x"3c032c22",
x"1c410c60",
x"fd8fedae",
x"ddcdcdec",
x"bd0bad2a",
x"9d498d68",
x"6eb67e97",
x"4ef45ed5",
x"2e323e13",
x"0e701e51",
x"efbeff9f",
x"cffcdfdd",
x"af3abf1b",
x"8f789f59",
x"81a99188",
x"a1ebb1ca",
x"c12dd10c",
x"e16ff14e",
x"00a11080",
x"20e330c2",
x"40255004",
x"60677046",
x"939883b9",
x"b3daa3fb",
x"d31cc33d",
x"f35ee37f",
x"129002b1",
x"32d222f3",
x"52144235",
x"72566277",
x"a5cbb5ea",
x"858995a8",
x"e54ff56e",
x"c50dd52c",
x"24c334e2",
x"048114a0",
x"64477466",
x"44055424",
x"b7faa7db",
x"97b88799",
x"f77ee75f",
x"d73cc71d",
x"36f226d3",
x"16b00691",
x"76766657",
x"56344615",
x"c96dd94c",
x"e92ff90e",
x"89e999c8",
x"a9abb98a",
x"48655844",
x"68277806",
x"08e118c0",
x"28a33882",
x"db5ccb7d",
x"fb1eeb3f",
x"9bd88bf9",
x"bb9aabbb",
x"5a544a75",
x"7a166a37",
x"1ad00af1",
x"3a922ab3",
x"ed0ffd2e",
x"cd4ddd6c",
x"ad8bbdaa",
x"8dc99de8",
x"6c077c26",
x"4c455c64",
x"2c833ca2",
x"0cc11ce0",
x"ff3eef1f",
x"df7ccf5d",
x"bfbaaf9b",
x"9ff88fd9",
x"7e366e17",
x"5e744e55",
x"3eb22e93",
x"1ef00ed1",
x"32313035",
x"00000000",
x"34333231",
x"00000000",
x"3437382d",
x"00000000",
x"3232312b",
x"00000000",
x"352e3533",
x"30303434",
x"00000000",
x"3332312e",
x"30303534",
x"00000000",
x"3031312d",
x"3030372e",
x"00000000",
x"362e302b",
x"30303434",
x"00000000",
x"30352e35",
x"332b6530",
x"00000000",
x"32312e2d",
x"322d6533",
x"00000000",
x"6537382d",
x"3233382b",
x"00000000",
x"362e302b",
x"32312d65",
x"00000000",
x"332e3054",
x"46312d65",
x"00000000",
x"542e542d",
x"71542b2b",
x"00000000",
x"2e335431",
x"7a346534",
x"00000000",
x"302e3433",
x"5e542d65",
x"00000000",
x"0000aed2",
x"0000b0b4",
x"0000af3e",
x"0000b020",
x"0000af92",
x"0000afd4",
x"0000b060",
x"0000b094",
x"0000b15e",
x"0000b120",
x"0000b12e",
x"0000b138",
x"0000b146",
x"0000b154",
x"ce221101",
x"26231000",
x"0793fea4",
x"439ce000",
x"4472853e",
x"80826105",
x"c6221141",
x"07930800",
x"4798e000",
x"8ff967a1",
x"4785c399",
x"4781a011",
x"4432853e",
x"80820141",
x"c6061141",
x"0800c422",
x"87aa3fe1",
x"40b2853e",
x"01414422",
x"71798082",
x"1800d622",
x"879377fd",
x"43dc4007",
x"fef42623",
x"879377fd",
x"439c4007",
x"fef42423",
x"879377fd",
x"43dc4007",
x"fef42223",
x"fec42703",
x"fe442783",
x"00f70363",
x"0001bfc1",
x"fe842783",
x"fcf42c23",
x"fe442783",
x"fcf42e23",
x"fd842703",
x"fdc42783",
x"85be853a",
x"61455432",
x"71798082",
x"1800d622",
x"fca42c23",
x"fcb42e23",
x"fd842703",
x"fdc42783",
x"fee42423",
x"fef42623",
x"879377fd",
x"577d4007",
x"77fdc798",
x"40078793",
x"fec42703",
x"77fdc7d8",
x"40078793",
x"fe842703",
x"0001c798",
x"54320001",
x"80826145",
x"ce221101",
x"77fd1000",
x"40078793",
x"2423479c",
x"77fdfef4",
x"40078793",
x"262347dc",
x"2703fef4",
x"2783fe84",
x"853afec4",
x"447285be",
x"80826105",
x"c6061141",
x"0800c422",
x"872a37e1",
x"853a87ae",
x"40b285be",
x"01414422",
x"11018082",
x"cc22ce06",
x"24231000",
x"2623fea4",
x"2503feb4",
x"2583fe84",
x"3f91fec4",
x"40f20001",
x"61054462",
x"11418082",
x"c422c606",
x"35d50800",
x"87ae872a",
x"85be853a",
x"442240b2",
x"80820141",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"00013057",
x"61054472",
x"11018082",
x"1000ce22",
x"342027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce221101",
x"27f31000",
x"26233420",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"feb42423",
x"fec42703",
x"f46347bd",
x"478500e7",
x"07b7a839",
x"87138000",
x"27830987",
x"078afec4",
x"270397ba",
x"c398fe84",
x"0000100f",
x"853e4781",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"feb42423",
x"fec42703",
x"f46347bd",
x"478500e7",
x"8713a829",
x"27838701",
x"078afec4",
x"270397ba",
x"c398fe84",
x"0000100f",
x"853e4781",
x"61054472",
x"71798082",
x"d422d606",
x"2e231800",
x"2783fca4",
x"9bf1fdc4",
x"fef42623",
x"fec42503",
x"00013f31",
x"542250b2",
x"80826145",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"ce86711d",
x"ca9acc96",
x"c6a2c89e",
x"c2aec4aa",
x"de36c0b2",
x"da3edc3a",
x"d646d842",
x"d276d472",
x"ce7ed07a",
x"35f11080",
x"faa42623",
x"fac42783",
x"242383fd",
x"2783faf4",
x"f793fac4",
x"22233ff7",
x"2703faf4",
x"4785fa84",
x"00f71d63",
x"800007b7",
x"09878713",
x"fa442783",
x"97ba078a",
x"9782439c",
x"8713a819",
x"27838701",
x"078afa44",
x"439c97ba",
x"fa442503",
x"00019782",
x"42e640f6",
x"43c64356",
x"45264436",
x"46064596",
x"576256f2",
x"584257d2",
x"5e2258b2",
x"5f025e92",
x"61254ff2",
x"30200073",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"ce061101",
x"1000cc22",
x"fe042623",
x"8713a005",
x"27838701",
x"078afec4",
x"672197ba",
x"16470713",
x"2783c398",
x"0785fec4",
x"fef42623",
x"fec42703",
x"fee347bd",
x"67a1fce7",
x"70078513",
x"000135bd",
x"446240f2",
x"80826105",
x"c6061141",
x"0800c422",
x"00013f45",
x"442240b2",
x"80820141",
x"ce061101",
x"1000cc22",
x"fea42623",
x"feb42423",
x"fe842583",
x"fec42503",
x"87aa3b6d",
x"40f2853e",
x"61054462",
x"11018082",
x"cc22ce06",
x"26231000",
x"2423fea4",
x"2583feb4",
x"2503fe84",
x"3bd1fec4",
x"853e87aa",
x"446240f2",
x"80826105",
x"ce221101",
x"87aa1000",
x"fef407a3",
x"77fd0001",
x"50078793",
x"07b74398",
x"8ff90020",
x"77fdfbed",
x"50078793",
x"fef44703",
x"0001c3d8",
x"61054472",
x"71798082",
x"d422d606",
x"2e231800",
x"2c23fca4",
x"20c1fcb4",
x"cbcd87aa",
x"fe042623",
x"fe042423",
x"879377fd",
x"a0235007",
x"27830007",
x"0786fd84",
x"fdc42703",
x"02f757b3",
x"fef42423",
x"2703a81d",
x"4789fec4",
x"00f70763",
x"fec42703",
x"18634791",
x"278300f7",
x"838dfe84",
x"fef42423",
x"2783a031",
x"8385fe84",
x"fef42423",
x"fec42783",
x"26230785",
x"2703fef4",
x"0793fe84",
x"e2e33fe0",
x"2223fce7",
x"2783fe04",
x"e793fe44",
x"22230017",
x"2783fef4",
x"078efec4",
x"27038be1",
x"8fd9fe44",
x"fef42223",
x"fe842783",
x"971317fd",
x"67c10067",
x"8ff917fd",
x"fe442703",
x"22238fd9",
x"77fdfef4",
x"50078793",
x"fe442703",
x"a011c398",
x"50b20001",
x"61455422",
x"11018082",
x"1000ce22",
x"fe042623",
x"e0000793",
x"07b74798",
x"8ff90002",
x"4785c781",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce061101",
x"1000cc22",
x"fea42623",
x"feb42423",
x"fe842583",
x"fec42503",
x"000135fd",
x"446240f2",
x"80826105",
x"ce061101",
x"1000cc22",
x"07a387aa",
x"4783fef4",
x"853efef4",
x"00013d71",
x"446240f2",
x"80826105",
x"d6227179",
x"d24ed44a",
x"2c231800",
x"2e23fca4",
x"2623fcb4",
x"2583fe04",
x"e581fdc4",
x"02000593",
x"4581a011",
x"feb42423",
x"fec42503",
x"fe842583",
x"262395aa",
x"2583feb4",
x"1581fe84",
x"0005c863",
x"fd842503",
x"00b51eb3",
x"a8154e01",
x"fd842583",
x"0015d513",
x"258342fd",
x"85b3fe84",
x"55b340b2",
x"250300b5",
x"2283fe84",
x"9eb3fdc4",
x"eeb300a2",
x"258301d5",
x"2503fe84",
x"1e33fd84",
x"2c2300b5",
x"2e23fdc4",
x"2503fdd4",
x"65c1fdc4",
x"00b57463",
x"a01145c1",
x"24234581",
x"2503feb4",
x"2583fec4",
x"95aafe84",
x"feb42623",
x"fe842583",
x"c8631581",
x"25030005",
x"13b3fd84",
x"430100b5",
x"2583a815",
x"d513fd84",
x"4e7d0015",
x"fe842583",
x"40be05b3",
x"00b555b3",
x"fe842503",
x"fdc42e03",
x"00ae13b3",
x"0075e3b3",
x"fe842583",
x"fd842503",
x"00b51333",
x"fc642c23",
x"fc742e23",
x"fdc42503",
x"010005b7",
x"00b57463",
x"a01145a1",
x"24234581",
x"2503feb4",
x"2583fec4",
x"95aafe84",
x"feb42623",
x"fe842583",
x"c8631581",
x"25030005",
x"18b3fd84",
x"480100b5",
x"2583a815",
x"d513fd84",
x"437d0015",
x"fe842583",
x"40b305b3",
x"00b555b3",
x"fe842503",
x"fdc42303",
x"00a318b3",
x"0115e8b3",
x"fe842583",
x"fd842503",
x"00b51833",
x"fd042c23",
x"fd142e23",
x"fdc42503",
x"100005b7",
x"00b57463",
x"a0114591",
x"24234581",
x"2503feb4",
x"2583fec4",
x"95aafe84",
x"feb42623",
x"fe842583",
x"c8631581",
x"25030005",
x"16b3fd84",
x"460100b5",
x"2583a80d",
x"d513fd84",
x"487d0015",
x"fe842583",
x"40b805b3",
x"00b555b3",
x"fe842503",
x"fdc42803",
x"00a816b3",
x"25838ecd",
x"2503fe84",
x"1633fd84",
x"2c2300b5",
x"2e23fcc4",
x"2603fcd4",
x"06b7fdc4",
x"74634000",
x"468900d6",
x"4681a011",
x"fed42423",
x"fec42603",
x"fe842683",
x"262396b2",
x"2683fed4",
x"1681fe84",
x"0006c863",
x"fd842603",
x"00d617b3",
x"a80d4701",
x"fd842683",
x"0016d613",
x"268345fd",
x"86b3fe84",
x"56b340d5",
x"260300d6",
x"2583fe84",
x"97b3fdc4",
x"8fd500c5",
x"fe842683",
x"fd842603",
x"00d61733",
x"fce42c23",
x"fcf42e23",
x"fd842703",
x"fdc42783",
x"fff74f13",
x"fff7cf93",
x"01ffd913",
x"77934981",
x"873e0ff9",
x"fec42783",
x"853e97ba",
x"59225432",
x"61455992",
x"71718082",
x"d522d706",
x"d14ad326",
x"cd52cf4e",
x"c95acb56",
x"c562c75e",
x"c16ac366",
x"1900deee",
x"f8a42c23",
x"f8b42e23",
x"f8c42823",
x"f8d42a23",
x"f8e42623",
x"f9442703",
x"f9c42783",
x"00e7ee63",
x"f9442703",
x"f9c42783",
x"02f71a63",
x"f9042703",
x"f9842783",
x"02e7f463",
x"f8c42783",
x"2683cb89",
x"2703f8c4",
x"2783f984",
x"c298f9c4",
x"4781c2dc",
x"20234801",
x"2223f8f4",
x"a681f904",
x"f9042703",
x"f9442783",
x"2783e3f9",
x"2703f904",
x"8fd9f944",
x"03a3e795",
x"4783fa04",
x"f793fa74",
x"873e0ff7",
x"078587ba",
x"0037b793",
x"0ff7f793",
x"87bac399",
x"4781a011",
x"0ff7f793",
x"faf403a3",
x"f9042703",
x"17634785",
x"278302f7",
x"e39df944",
x"f8c42783",
x"2783c799",
x"4681f8c4",
x"c3944701",
x"2783c3d8",
x"2803f984",
x"2023f9c4",
x"2223f8f4",
x"a4f1f904",
x"f9842703",
x"f9c42783",
x"2783eba9",
x"c78df8c4",
x"f9842703",
x"f9c42783",
x"270386ba",
x"2783f904",
x"87baf944",
x"02f6f7b3",
x"4881883e",
x"f8c42783",
x"0107a023",
x"0117a223",
x"f9842703",
x"f9c42783",
x"270386ba",
x"2783f904",
x"87baf944",
x"02f6d7b3",
x"f8f42023",
x"f8042223",
x"2503ac8d",
x"2583f904",
x"390df944",
x"f49387aa",
x"25030ff7",
x"2583f984",
x"310df9c4",
x"f79387aa",
x"87b30ff7",
x"f79340f4",
x"07850ff7",
x"faf40fa3",
x"fbf44783",
x"fe078713",
x"00074863",
x"f9c42783",
x"00e7da33",
x"a01d4a81",
x"f9c42703",
x"00171693",
x"8f1d477d",
x"00e69733",
x"f9842683",
x"00f6da33",
x"01476a33",
x"f9c42703",
x"00f75ab3",
x"fb442823",
x"fb542a23",
x"fbf44783",
x"04000713",
x"40f707b3",
x"fe078713",
x"00074863",
x"f9842783",
x"00e799b3",
x"a01d4901",
x"f9842703",
x"00175693",
x"8f1d477d",
x"00e6d733",
x"f9c42683",
x"00f699b3",
x"013769b3",
x"f9842703",
x"00f71933",
x"f9242c23",
x"f9342e23",
x"48014781",
x"faf42423",
x"fb042623",
x"2783aa1d",
x"83fdfb04",
x"fb442703",
x"00171c93",
x"0197ecb3",
x"fb042783",
x"00179c13",
x"f9c42783",
x"2c2383fd",
x"2e23f6f4",
x"2683f604",
x"2703f784",
x"87b6f7c4",
x"00fc67b3",
x"faf42823",
x"e7b387ba",
x"2a2300fc",
x"2783faf4",
x"83fdf984",
x"f9c42703",
x"00171d93",
x"01b7edb3",
x"f9842783",
x"00179d13",
x"fa842783",
x"28238b85",
x"2783f6f4",
x"8b81fac4",
x"f6f42a23",
x"f7042683",
x"f7442703",
x"67b387b6",
x"2c2300fd",
x"87baf8f4",
x"00fde7b3",
x"f8f42e23",
x"f9042703",
x"f9442783",
x"fb042503",
x"fb442583",
x"40a70633",
x"38338832",
x"86b30107",
x"87b340b7",
x"86be4106",
x"55fd557d",
x"00a60733",
x"3833883a",
x"87b300c8",
x"06b300b6",
x"87b600f8",
x"41f7d693",
x"f6d42423",
x"262387fd",
x"2783f6f4",
x"2803f684",
x"2423f6c4",
x"2623faf4",
x"2703fb04",
x"2783f904",
x"8ff9fa84",
x"f6f42023",
x"f9442703",
x"fac42783",
x"22238ff9",
x"2603f6f4",
x"2683fb04",
x"2803fb44",
x"2883f604",
x"85c2f644",
x"40b60733",
x"35b385ba",
x"854600b6",
x"40a687b3",
x"40b786b3",
x"282387b6",
x"2a23fae4",
x"4783faf4",
x"8713fbf4",
x"0fa3fff7",
x"90e3fae4",
x"2783ec07",
x"cb89f8c4",
x"f8c42683",
x"fb042703",
x"fb442783",
x"c2dcc298",
x"f9842783",
x"270383fd",
x"1b93f9c4",
x"ebb30017",
x"27830177",
x"9b13f984",
x"27830017",
x"8b85fa84",
x"f4f42c23",
x"fac42783",
x"2e238b81",
x"2683f4f4",
x"2703f584",
x"87b6f5c4",
x"00fb67b3",
x"f8f42023",
x"e7b387ba",
x"222300fb",
x"2703f8f4",
x"2783f804",
x"853af844",
x"50ba85be",
x"549a542a",
x"49fa590a",
x"4ada4a6a",
x"4bba4b4a",
x"4c9a4c2a",
x"5df64d0a",
x"8082614d",
x"ce061101",
x"1000cc22",
x"fea42423",
x"feb42623",
x"fec42023",
x"fed42223",
x"26034701",
x"2683fe04",
x"2503fe44",
x"2583fe84",
x"3ed5fec4",
x"87ae872a",
x"85be853a",
x"446240f2",
x"80826105",
x"d6227179",
x"2e231800",
x"2c23fca4",
x"57fdfcb4",
x"fef41723",
x"fe042423",
x"2783a8a9",
x"2703fe84",
x"97bafdc4",
x"0007c703",
x"fee45783",
x"07c283a1",
x"f79383c1",
x"8fb90ff7",
x"fef403a3",
x"fe744783",
x"07136721",
x"07861747",
x"d78397ba",
x"97130007",
x"87410107",
x"fee41783",
x"07c207a2",
x"8fb987c1",
x"87c107c2",
x"fef41723",
x"fe842783",
x"24230785",
x"2703fef4",
x"2783fe84",
x"40e3fd84",
x"5783faf7",
x"853efee4",
x"61455432",
x"71798082",
x"d422d606",
x"2e231800",
x"87aefca4",
x"fcc42a23",
x"fcf40da3",
x"fdc42783",
x"faa00713",
x"00e78023",
x"fdc42783",
x"fdb44703",
x"00e780a3",
x"fdc42783",
x"00078123",
x"0793a82d",
x"85befef4",
x"fd442503",
x"87aa2c49",
x"2783c78d",
x"c783fdc4",
x"87130027",
x"76930017",
x"27030ff7",
x"0123fdc4",
x"86be00d7",
x"fef44703",
x"fdc42783",
x"81a397b6",
x"250300e7",
x"2a91fd44",
x"c79387aa",
x"f7930017",
x"cb890ff7",
x"fdc42783",
x"0027c703",
x"0ff00793",
x"faf715e3",
x"fdc42783",
x"00378713",
x"fdc42783",
x"0027c783",
x"853a85be",
x"87aa3dc1",
x"2783873e",
x"9123fdc4",
x"278310e7",
x"0713fdc4",
x"82230550",
x"000110e7",
x"542250b2",
x"80826145",
x"d6067179",
x"1800d422",
x"fca42e23",
x"fdc42783",
x"0007c783",
x"f0ef853e",
x"2783fdaf",
x"c783fdc4",
x"853e0017",
x"fccff0ef",
x"fdc42783",
x"0027c783",
x"f0ef853e",
x"2623fbef",
x"a005fe04",
x"fdc42703",
x"fec42783",
x"c78397ba",
x"853e0037",
x"fa4ff0ef",
x"fec42783",
x"26230785",
x"2783fef4",
x"c783fdc4",
x"873e0027",
x"fec42783",
x"fce7eae3",
x"fdc42783",
x"1027d783",
x"07c283a1",
x"f79383c1",
x"853e0ff7",
x"f70ff0ef",
x"fdc42783",
x"1027d783",
x"0ff7f793",
x"f0ef853e",
x"2783f5ef",
x"c783fdc4",
x"853e1047",
x"f50ff0ef",
x"50b20001",
x"61455422",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"10079023",
x"fec42783",
x"10079123",
x"fec42783",
x"10079223",
x"44720001",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"d783fec4",
x"87931047",
x"b793f007",
x"f7930017",
x"853e0ff7",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"1047d783",
x"0017b793",
x"0ff7f793",
x"4472853e",
x"80826105",
x"d6067179",
x"1800d422",
x"fca42e23",
x"fcb42c23",
x"fe042623",
x"2783a82d",
x"078efec4",
x"fd842703",
x"00f757b3",
x"fef405a3",
x"feb44783",
x"250385be",
x"280dfdc4",
x"c79387aa",
x"f7930017",
x"c3990ff7",
x"a8214781",
x"fec42783",
x"26230785",
x"2703fef4",
x"478dfec4",
x"fce7d1e3",
x"853e4785",
x"542250b2",
x"80826145",
x"ce061101",
x"1000cc22",
x"fea42623",
x"05a387ae",
x"2503fef4",
x"3f3dfec4",
x"c39987aa",
x"a8b94781",
x"fec42783",
x"1027d783",
x"2783873e",
x"97bafec4",
x"feb44703",
x"00e78023",
x"fec42783",
x"1027d783",
x"00178713",
x"41f75793",
x"973e83e1",
x"0ff77713",
x"40f707b3",
x"01079713",
x"27838341",
x"9123fec4",
x"278310e7",
x"d783fec4",
x"07851047",
x"01079713",
x"27838341",
x"9223fec4",
x"478510e7",
x"40f2853e",
x"61054462",
x"11018082",
x"cc22ce06",
x"26231000",
x"2423fea4",
x"2503feb4",
x"35c5fec4",
x"c39987aa",
x"a08d4781",
x"fec42783",
x"1007d783",
x"2783873e",
x"97bafec4",
x"0007c703",
x"fe842783",
x"00e78023",
x"fec42783",
x"1007d783",
x"00178713",
x"41f75793",
x"973e83e1",
x"0ff77713",
x"40f707b3",
x"01079713",
x"27838341",
x"9023fec4",
x"278310e7",
x"d783fec4",
x"17fd1047",
x"01079713",
x"27838341",
x"9223fec4",
x"478510e7",
x"40f2853e",
x"61054462",
x"11018082",
x"1000ce22",
x"fea42623",
x"feb42423",
x"fe842783",
x"00079703",
x"fec42783",
x"00e79023",
x"fe842783",
x"00279703",
x"fec42783",
x"00e79123",
x"44720001",
x"80826105",
x"c686715d",
x"0880c4a2",
x"faa42e23",
x"fab42c23",
x"1b2387b2",
x"47d1faf4",
x"fef42223",
x"fbc42703",
x"fe442783",
x"02f757b3",
x"202317f9",
x"2703fef4",
x"2783fb84",
x"078efe04",
x"2e2397ba",
x"2783fcf4",
x"2423fdc4",
x"2703fcf4",
x"2783fc84",
x"078afe04",
x"2c2397ba",
x"2783fcf4",
x"2a23fb84",
x"2783fcf4",
x"a023fd44",
x"27030007",
x"2783fc84",
x"c3d8fd44",
x"fd442783",
x"912343dc",
x"27830007",
x"43dcfd44",
x"07137761",
x"90230807",
x"278300e7",
x"07a1fb84",
x"faf42c23",
x"fc842783",
x"24230791",
x"77e1fcf4",
x"fff7c793",
x"fcf41323",
x"122357fd",
x"0693fcf4",
x"0613fc84",
x"0593fb84",
x"2783fc44",
x"2703fd84",
x"2503fdc4",
x"2a91fd44",
x"fe042623",
x"2783a8ad",
x"9713fec4",
x"83410107",
x"fb645783",
x"07c28fb9",
x"8bbd83c1",
x"fcf41823",
x"fd045783",
x"9713078e",
x"83410107",
x"fec42783",
x"83c107c2",
x"07c28b9d",
x"8fd983c1",
x"fcf41723",
x"fce41783",
x"971307a2",
x"87410107",
x"fce41783",
x"07c28fd9",
x"122387c1",
x"0693fcf4",
x"0613fc84",
x"0593fb84",
x"2783fc44",
x"2703fd84",
x"2503fdc4",
x"20c5fd44",
x"fec42783",
x"26230785",
x"2703fef4",
x"2783fec4",
x"60e3fe04",
x"2783f8f7",
x"439cfd44",
x"fef42423",
x"26234785",
x"a841fef4",
x"fe042703",
x"57b34795",
x"270302f7",
x"7063fec4",
x"278302f7",
x"8713fec4",
x"26230017",
x"2703fee4",
x"4358fe84",
x"87c107c2",
x"00f71123",
x"2783a8a1",
x"8713fec4",
x"26230017",
x"9713fee4",
x"83410107",
x"fb645783",
x"19238fb9",
x"2783fcf4",
x"07c2fec4",
x"07a283c1",
x"83c107c2",
x"7007f793",
x"83c107c2",
x"fd245703",
x"07c28fd9",
x"969383c1",
x"86c10107",
x"fe842783",
x"671143dc",
x"8f75177d",
x"87410742",
x"00e79123",
x"fe842783",
x"2423439c",
x"2783fef4",
x"439cfe84",
x"4601f7b5",
x"5b400593",
x"fd442503",
x"cf3f60ef",
x"fca42a23",
x"fd442783",
x"40b6853e",
x"61614426",
x"71398082",
x"dc22de06",
x"2e230080",
x"2c23fca4",
x"2a23fcb4",
x"2823fcc4",
x"2623fcd4",
x"2423fce4",
x"2783fcf4",
x"439cfd44",
x"270307a1",
x"e463fcc4",
x"478100e7",
x"2783a895",
x"439cfd04",
x"27030791",
x"e463fc84",
x"478100e7",
x"2783a085",
x"439cfd44",
x"fef42623",
x"fd442783",
x"8713439c",
x"27830087",
x"c398fd44",
x"fdc42783",
x"27834398",
x"c398fec4",
x"fdc42783",
x"fec42703",
x"2783c398",
x"4398fd04",
x"fec42783",
x"2783c3d8",
x"439cfd04",
x"00478713",
x"fd042783",
x"2783c398",
x"43dcfec4",
x"fd842583",
x"3b01853e",
x"fec42783",
x"50f2853e",
x"61215462",
x"71398082",
x"dc22de06",
x"0080da26",
x"fca42623",
x"fcb42423",
x"fe041623",
x"fe041523",
x"142357fd",
x"1323fef4",
x"1b23fe04",
x"4505fc04",
x"13d010ef",
x"971387aa",
x"87410107",
x"fcc42783",
x"00e79023",
x"10ef4509",
x"87aa1270",
x"01079713",
x"27838741",
x"9123fcc4",
x"450d00e7",
x"111010ef",
x"971387aa",
x"87410107",
x"fcc42783",
x"00e79223",
x"10ef4511",
x"87aa0fb0",
x"2783873e",
x"cfd8fcc4",
x"10ef4515",
x"87aa0eb0",
x"2783873e",
x"d398fcc4",
x"fcc42783",
x"e789539c",
x"fcc42783",
x"d398471d",
x"fcc42783",
x"00079783",
x"2783eb8d",
x"9783fcc4",
x"e7850027",
x"fcc42783",
x"00479783",
x"2783ef99",
x"9023fcc4",
x"27830007",
x"9123fcc4",
x"27830007",
x"0713fcc4",
x"92230660",
x"278300e7",
x"9703fcc4",
x"47850007",
x"04f71063",
x"fcc42783",
x"00279783",
x"2783eb95",
x"9783fcc4",
x"e78d0047",
x"fcc42783",
x"0713670d",
x"90234157",
x"278300e7",
x"670dfcc4",
x"41570713",
x"00e79123",
x"fcc42783",
x"06600713",
x"00e79223",
x"fcc42783",
x"80000737",
x"11870713",
x"2783c798",
x"0713fcc4",
x"cf987d00",
x"fcc42783",
x"04079023",
x"fe041723",
x"5783a035",
x"4705fee4",
x"00f717b3",
x"2783873e",
x"539cfcc4",
x"c7918ff9",
x"fea45783",
x"15230785",
x"5783fef4",
x"0785fee4",
x"fef41723",
x"fee45703",
x"f8e34789",
x"1723fce7",
x"a081fe04",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafcc4",
x"56834f90",
x"5703fea4",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fcc42783",
x"573397ba",
x"cf9802d6",
x"fee45783",
x"17230785",
x"5783fef4",
x"dfddfee4",
x"fe041723",
x"5783a071",
x"4705fee4",
x"00f717b3",
x"2783873e",
x"539cfcc4",
x"c7b58ff9",
x"fe042023",
x"2703a899",
x"87bafe04",
x"97ba0792",
x"873e078a",
x"fcc42783",
x"478c97ba",
x"fcc42783",
x"57834f98",
x"0633fec4",
x"270302f7",
x"87bafe04",
x"97ba0792",
x"873e078a",
x"fcc42783",
x"00e786b3",
x"fee45783",
x"87330785",
x"078a00c5",
x"c79897b6",
x"fe042783",
x"20230785",
x"2783fef4",
x"d7c5fe04",
x"fec45783",
x"16230785",
x"5783fef4",
x"0785fee4",
x"fef41723",
x"fee45703",
x"f8e34789",
x"1723f6e7",
x"aaa9fe04",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafcc4",
x"8b85539c",
x"2783cbb1",
x"4f94fcc4",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafcc4",
x"570347cc",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fcc42783",
x"960397ba",
x"57030007",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fcc42783",
x"00e784b3",
x"34bd8536",
x"d0dc87aa",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafcc4",
x"8b89539c",
x"2783cbb5",
x"4f88fcc4",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafcc4",
x"57034b8c",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fcc42783",
x"978397ba",
x"86be0007",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafcc4",
x"00279783",
x"e63307c2",
x"570300f6",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fcc42783",
x"879397ba",
x"86be0287",
x"dd1f60ef",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafcc4",
x"8b91539c",
x"2783cf9d",
x"4f94fcc4",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafcc4",
x"00079583",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafcc4",
x"863e4bdc",
x"10ef8536",
x"57831180",
x"0785fee4",
x"fef41723",
x"fee45783",
x"ea0782e3",
x"fcc42783",
x"e3d14fdc",
x"fc042e23",
x"fcc42783",
x"cfd84705",
x"2783a081",
x"4fd8fcc4",
x"078a87ba",
x"078697ba",
x"2783873e",
x"cfd8fcc4",
x"64d000ef",
x"fcc42503",
x"c59f60ef",
x"665000ef",
x"685000ef",
x"87ae872a",
x"fc842603",
x"85be853a",
x"6b9000ef",
x"fca42e23",
x"fdc42783",
x"2783dfdd",
x"2c23fdc4",
x"2783fcf4",
x"e781fd84",
x"2c234785",
x"2783fcf4",
x"4fd8fcc4",
x"278346a9",
x"d7b3fd84",
x"078502f6",
x"02f70733",
x"fcc42783",
x"00efcfd8",
x"25035ef0",
x"60effcc4",
x"00efbfbf",
x"27836070",
x"9783fcc4",
x"57030007",
x"85bafd64",
x"70ef853e",
x"87aa9d4f",
x"fcf41b23",
x"fcc42783",
x"00279783",
x"fd645703",
x"853e85ba",
x"9baf70ef",
x"1b2387aa",
x"2783fcf4",
x"9783fcc4",
x"57030047",
x"85bafd64",
x"70ef853e",
x"87aa9a0f",
x"fcf41b23",
x"fcc42783",
x"07c24f9c",
x"570387c1",
x"85bafd64",
x"70ef853e",
x"87aa984f",
x"fcf41b23",
x"fd645783",
x"0713673d",
x"81639f57",
x"673d06e7",
x"9f570713",
x"06f74463",
x"07136725",
x"8c63a027",
x"672502e7",
x"a0270713",
x"04f74a63",
x"07136721",
x"8563b057",
x"672102e7",
x"b0570713",
x"04f74063",
x"07136709",
x"87638f27",
x"671502e7",
x"eaf70713",
x"00e78a63",
x"1423a025",
x"a02dfe04",
x"14234785",
x"a00dfef4",
x"14234789",
x"a829fef4",
x"1423478d",
x"a809fef4",
x"14234791",
x"a029fef4",
x"132357fd",
x"0001fef4",
x"fe841783",
x"1c07c263",
x"fe041723",
x"5703a275",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fcc42783",
x"902397ba",
x"57030407",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fcc42783",
x"539c97ba",
x"cfb18b85",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafcc4",
x"03a7d703",
x"fe841783",
x"800006b7",
x"00068693",
x"97b60786",
x"0007d783",
x"02f70763",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafcc4",
x"04079703",
x"83410742",
x"07420705",
x"07428341",
x"90238741",
x"570304e7",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fcc42783",
x"539c97ba",
x"cfb18b89",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafcc4",
x"03c7d703",
x"fe841783",
x"800006b7",
x"00c68693",
x"97b60786",
x"0007d783",
x"02f70763",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafcc4",
x"04079703",
x"83410742",
x"07420705",
x"07428341",
x"90238741",
x"570304e7",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fcc42783",
x"539c97ba",
x"cfb18b91",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafcc4",
x"03e7d703",
x"fe841783",
x"800006b7",
x"01868693",
x"97b60786",
x"0007d783",
x"02f70763",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafcc4",
x"04079703",
x"83410742",
x"07420705",
x"07428341",
x"90238741",
x"570304e7",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fcc42783",
x"978397ba",
x"97130407",
x"83410107",
x"fe645783",
x"07c297ba",
x"132383c1",
x"5783fef4",
x"0785fee4",
x"fef41723",
x"fee45703",
x"800007b7",
x"0707a783",
x"e4f765e3",
x"fe641783",
x"50f2853e",
x"54d25462",
x"80826121",
x"de067139",
x"0080dc22",
x"fca42e23",
x"fcb42c23",
x"fcc42a23",
x"fcd42823",
x"172387ba",
x"1723fcf4",
x"5783fe04",
x"873efce4",
x"8fd977fd",
x"fef41623",
x"fce41783",
x"2583863e",
x"2503fd44",
x"2469fdc4",
x"fce41783",
x"260386be",
x"2583fd44",
x"2503fd84",
x"2ae1fdc4",
x"fec41783",
x"2583863e",
x"2503fd84",
x"20edfdc4",
x"873e87aa",
x"fee45783",
x"853a85be",
x"eaff60ef",
x"172387aa",
x"2683fef4",
x"2603fd04",
x"2583fd44",
x"2503fd84",
x"24e5fdc4",
x"fec41783",
x"2583863e",
x"2503fd84",
x"284dfdc4",
x"873e87aa",
x"fee45783",
x"853a85be",
x"e77f60ef",
x"172387aa",
x"2683fef4",
x"2603fd04",
x"2583fd44",
x"2503fd84",
x"26adfdc4",
x"fec41783",
x"2583863e",
x"2503fd84",
x"28adfdc4",
x"873e87aa",
x"fee45783",
x"853a85be",
x"e3ff60ef",
x"172387aa",
x"2683fef4",
x"2603fd04",
x"2583fd44",
x"2503fd84",
x"2181fdc4",
x"fec41783",
x"2583863e",
x"2503fd84",
x"2089fdc4",
x"873e87aa",
x"fee45783",
x"853a85be",
x"e07f60ef",
x"172387aa",
x"5783fef4",
x"07b3fce4",
x"07c240f0",
x"07c283c1",
x"863e87c1",
x"fd442583",
x"fdc42503",
x"17832271",
x"853efee4",
x"546250f2",
x"80826121",
x"de227139",
x"26230080",
x"2423fca4",
x"87b2fcb4",
x"fcf41323",
x"fe042623",
x"fe042423",
x"fc042c23",
x"fe041323",
x"fe042023",
x"2e23a879",
x"a049fc04",
x"fe042703",
x"fcc42783",
x"02f70733",
x"fdc42783",
x"078a97ba",
x"fc842703",
x"439c97ba",
x"fcf42c23",
x"fec42703",
x"fd842783",
x"262397ba",
x"1783fef4",
x"2703fc64",
x"dc63fec4",
x"578300e7",
x"07a9fe64",
x"83c107c2",
x"fef41323",
x"fe042623",
x"2703a00d",
x"2783fd84",
x"a7b3fe84",
x"f79300e7",
x"873e0ff7",
x"fe645783",
x"07c297ba",
x"132383c1",
x"2783fef4",
x"2423fd84",
x"2783fef4",
x"0785fdc4",
x"fcf42e23",
x"fdc42703",
x"fcc42783",
x"f6f76ce3",
x"fe042783",
x"20230785",
x"2703fef4",
x"2783fe04",
x"6ee3fcc4",
x"1783f4f7",
x"853efe64",
x"61215472",
x"71798082",
x"1800d622",
x"fca42e23",
x"fcb42c23",
x"fcc42a23",
x"192387b6",
x"2623fcf4",
x"a0b5fe04",
x"fe042423",
x"2703a881",
x"2783fec4",
x"0733fdc4",
x"278302f7",
x"97bafe84",
x"27030786",
x"97bafd44",
x"00079783",
x"1703863e",
x"2683fd24",
x"2783fec4",
x"86b3fdc4",
x"278302f6",
x"97b6fe84",
x"2683078a",
x"97b6fd84",
x"02e60733",
x"2783c398",
x"0785fe84",
x"fef42423",
x"fe842703",
x"fdc42783",
x"faf765e3",
x"fec42783",
x"26230785",
x"2703fef4",
x"2783fec4",
x"67e3fdc4",
x"0001f8f7",
x"54320001",
x"80826145",
x"d6227179",
x"2e231800",
x"2c23fca4",
x"87b2fcb4",
x"fcf41b23",
x"fe042623",
x"2423a8b5",
x"a085fe04",
x"fec42703",
x"fdc42783",
x"02f70733",
x"fe842783",
x"078697ba",
x"fd842703",
x"978397ba",
x"97130007",
x"83410107",
x"fd645783",
x"969397ba",
x"82c10107",
x"fec42703",
x"fdc42783",
x"02f70733",
x"fe842783",
x"078697ba",
x"fd842703",
x"971397ba",
x"87410106",
x"00e79023",
x"fe842783",
x"24230785",
x"2703fef4",
x"2783fe84",
x"6de3fdc4",
x"2783f8f7",
x"0785fec4",
x"fef42623",
x"fec42703",
x"fdc42783",
x"f6f76fe3",
x"00010001",
x"61455432",
x"71798082",
x"1800d622",
x"fca42e23",
x"fcb42c23",
x"fcc42a23",
x"fcd42823",
x"fe042623",
x"2783a069",
x"078afec4",
x"fd842703",
x"a02397ba",
x"24230007",
x"a8b9fe04",
x"fec42783",
x"2703078a",
x"97bafd84",
x"27034394",
x"2783fec4",
x"0733fdc4",
x"278302f7",
x"97bafe84",
x"27030786",
x"97bafd44",
x"00079783",
x"2783863e",
x"0786fe84",
x"fd042703",
x"978397ba",
x"07330007",
x"278302f6",
x"078afec4",
x"fd842603",
x"973697b2",
x"2783c398",
x"0785fe84",
x"fef42423",
x"fe842703",
x"fdc42783",
x"f8f76ee3",
x"fec42783",
x"26230785",
x"2703fef4",
x"2783fec4",
x"68e3fdc4",
x"0001f6f7",
x"54320001",
x"80826145",
x"d6227179",
x"2e231800",
x"2c23fca4",
x"2a23fcb4",
x"2823fcc4",
x"2623fcd4",
x"a8f9fe04",
x"fe042423",
x"2703a0c9",
x"2783fec4",
x"0733fdc4",
x"278302f7",
x"97bafe84",
x"2703078a",
x"97bafd84",
x"0007a023",
x"fe042223",
x"2703a061",
x"2783fec4",
x"0733fdc4",
x"278302f7",
x"97bafe84",
x"2703078a",
x"97bafd84",
x"27034394",
x"2783fec4",
x"0733fdc4",
x"278302f7",
x"97bafe44",
x"27030786",
x"97bafd44",
x"00079783",
x"2703863e",
x"2783fe44",
x"0733fdc4",
x"278302f7",
x"97bafe84",
x"27030786",
x"97bafd04",
x"00079783",
x"02f60733",
x"fec42603",
x"fdc42783",
x"02f60633",
x"fe842783",
x"078a97b2",
x"fd842603",
x"973697b2",
x"2783c398",
x"0785fe44",
x"fef42223",
x"fe442703",
x"fdc42783",
x"f6f769e3",
x"fe842783",
x"24230785",
x"2703fef4",
x"2783fe84",
x"6ce3fdc4",
x"2783f2f7",
x"0785fec4",
x"fef42623",
x"fec42703",
x"fdc42783",
x"f0f76ee3",
x"00010001",
x"61455432",
x"71798082",
x"1800d622",
x"fca42e23",
x"fcb42c23",
x"fcc42a23",
x"fcd42823",
x"fe042623",
x"2423a8fd",
x"a0cdfe04",
x"fec42703",
x"fdc42783",
x"02f70733",
x"fe842783",
x"078a97ba",
x"fd842703",
x"a02397ba",
x"22230007",
x"a065fe04",
x"fec42703",
x"fdc42783",
x"02f70733",
x"fe442783",
x"078697ba",
x"fd442703",
x"978397ba",
x"86be0007",
x"fe442703",
x"fdc42783",
x"02f70733",
x"fe842783",
x"078697ba",
x"fd042703",
x"978397ba",
x"87b30007",
x"202302f6",
x"2703fef4",
x"2783fec4",
x"0733fdc4",
x"278302f7",
x"97bafe84",
x"2703078a",
x"97bafd84",
x"86be439c",
x"fe042783",
x"f7138789",
x"278300f7",
x"8795fe04",
x"07f7f793",
x"02f707b3",
x"270396be",
x"2783fec4",
x"0733fdc4",
x"278302f7",
x"97bafe84",
x"2703078a",
x"97bafd84",
x"c3988736",
x"fe442783",
x"22230785",
x"2703fef4",
x"2783fe44",
x"69e3fdc4",
x"2783f4f7",
x"0785fe84",
x"fef42423",
x"fe842703",
x"fdc42783",
x"f0f76ce3",
x"fec42783",
x"26230785",
x"2703fef4",
x"2783fec4",
x"6ee3fdc4",
x"0001eef7",
x"54320001",
x"80826145",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"00013207",
x"61054472",
x"11018082",
x"1000ce22",
x"b00027f3",
x"fef42623",
x"fec42783",
x"4681863e",
x"87b68732",
x"85be853a",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"b0079073",
x"44720001",
x"80826105",
x"ce221101",
x"27f31000",
x"2623b020",
x"2783fef4",
x"863efec4",
x"87324681",
x"853a87b6",
x"447285be",
x"80826105",
x"ce221101",
x"27f31000",
x"2623b030",
x"2783fef4",
x"863efec4",
x"87324681",
x"853a87b6",
x"447285be",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"0001b037",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"32379073",
x"44720001",
x"80826105",
x"ce221101",
x"27f31000",
x"2623c000",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"c80027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce221101",
x"27f31000",
x"2623b040",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"b0479073",
x"44720001",
x"80826105",
x"ce221101",
x"27f31000",
x"2623b050",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"b0579073",
x"44720001",
x"80826105",
x"ce221101",
x"27f31000",
x"2623b060",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"b0679073",
x"44720001",
x"80826105",
x"ce221101",
x"27f31000",
x"2623b070",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"b0779073",
x"44720001",
x"80826105",
x"ce221101",
x"27f31000",
x"2623b080",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"b0879073",
x"44720001",
x"80826105",
x"ce221101",
x"27f31000",
x"2623b090",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"b0979073",
x"44720001",
x"80826105",
x"ce221101",
x"27f31000",
x"2623b0a0",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"b0a79073",
x"44720001",
x"80826105",
x"ce221101",
x"27f31000",
x"2623b0b0",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"b0b79073",
x"44720001",
x"80826105",
x"ce221101",
x"27f31000",
x"2623b0c0",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"b0c79073",
x"44720001",
x"80826105",
x"ce221101",
x"27f31000",
x"2623b0d0",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"b0d79073",
x"44720001",
x"80826105",
x"ce221101",
x"27f31000",
x"2623b0e0",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"b0e79073",
x"44720001",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"00013247",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"32579073",
x"44720001",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"00013267",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"32779073",
x"44720001",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"00013287",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"32979073",
x"44720001",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"000132a7",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"32b79073",
x"44720001",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"000132c7",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"32d79073",
x"44720001",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"000132e7",
x"61054472",
x"71798082",
x"d422d606",
x"31511800",
x"fea42623",
x"24233195",
x"39a5fea4",
x"fea42223",
x"fec42703",
x"fe442783",
x"00f70363",
x"0001b7cd",
x"fe842783",
x"fcf42c23",
x"fe442783",
x"fcf42e23",
x"fd842703",
x"fdc42783",
x"85be853a",
x"542250b2",
x"80826145",
x"c6061141",
x"0800c422",
x"872a376d",
x"a02387ae",
x"a22382e1",
x"450182f1",
x"00013e25",
x"442240b2",
x"80820141",
x"c6061141",
x"0800c422",
x"360d557d",
x"872a3749",
x"a42387ae",
x"a62382e1",
x"000182f1",
x"442240b2",
x"80820141",
x"ce221101",
x"a6031000",
x"a6838281",
x"a50382c1",
x"a5838201",
x"07338241",
x"883a40a6",
x"01063833",
x"40b687b3",
x"410786b3",
x"242387b6",
x"2623fee4",
x"2703fef4",
x"2783fe84",
x"853afec4",
x"447285be",
x"80826105",
x"d6067179",
x"1800d422",
x"fca42c23",
x"fcb42e23",
x"fcc42a23",
x"fd442683",
x"47818736",
x"86be863a",
x"fd842503",
x"fdc42583",
x"df0fe0ef",
x"87ae872a",
x"fee42623",
x"fec42783",
x"50b2853e",
x"61455422",
x"11018082",
x"cc22ce06",
x"26231000",
x"2423fea4",
x"557dfeb4",
x"45013c85",
x"4501346d",
x"45213621",
x"45013e39",
x"45413649",
x"45013345",
x"0513367d",
x"3b450200",
x"3ee14501",
x"04000513",
x"450133c1",
x"05133109",
x"3bc10800",
x"31354501",
x"10000513",
x"450133c5",
x"05133999",
x"3bc52000",
x"31414501",
x"40000513",
x"45013501",
x"6785316d",
x"80078513",
x"45013539",
x"650539c9",
x"45013505",
x"650939fd",
x"45013d0d",
x"6511332d",
x"27833591",
x"4705fec4",
x"00e78023",
x"40f20001",
x"61054462",
x"71698082",
x"12112623",
x"12812423",
x"2e231a00",
x"2c23eca4",
x"2783ecb4",
x"8023edc4",
x"25830007",
x"8513ed84",
x"e0ef0801",
x"3ae1fc6f",
x"87ae872a",
x"85be87ba",
x"08018513",
x"fb4fe0ef",
x"872a3411",
x"87ba87ae",
x"851385be",
x"e0ef0801",
x"3c19fa2f",
x"87ae872a",
x"85be87ba",
x"08018513",
x"f90fe0ef",
x"87aa3c41",
x"851385be",
x"e0ef0801",
x"3c5df82f",
x"85be87aa",
x"08018513",
x"f74fe0ef",
x"87aa3cf1",
x"851385be",
x"e0ef0801",
x"3609f66f",
x"85be87aa",
x"08018513",
x"f58fe0ef",
x"87aa3625",
x"851385be",
x"e0ef0801",
x"36b9f4af",
x"85be87aa",
x"08018513",
x"f3cfe0ef",
x"87aa3e95",
x"851385be",
x"e0ef0801",
x"3e69f2ef",
x"85be87aa",
x"08018513",
x"f20fe0ef",
x"87aa36c1",
x"851385be",
x"e0ef0801",
x"36ddf12f",
x"85be87aa",
x"08018513",
x"f04fe0ef",
x"87aa3131",
x"851385be",
x"e0ef0801",
x"0713ef6f",
x"8613ee84",
x"45850801",
x"e0ef853a",
x"0793cfcf",
x"853eee84",
x"dbcfe0ef",
x"20830001",
x"240312c1",
x"61551281",
x"71798082",
x"1800d622",
x"fca42e23",
x"2a2387ae",
x"1d23fcc4",
x"2623fcf4",
x"2423fe04",
x"2023fe04",
x"2783fe04",
x"17fdfdc4",
x"fcf42e23",
x"fe042423",
x"2783a285",
x"c7a5fe84",
x"fe042223",
x"2703a03d",
x"2783fe04",
x"973efe44",
x"fec42683",
x"fe442783",
x"268397b6",
x"97b6fd44",
x"00074703",
x"00e78023",
x"fe442783",
x"22230785",
x"2703fef4",
x"2783fe44",
x"66e3fe84",
x"2703fcf7",
x"2783fec4",
x"97bafe44",
x"fd442703",
x"071397ba",
x"802302c0",
x"270300e7",
x"2783fe84",
x"97bafec4",
x"26230785",
x"1783fef4",
x"07c2fda4",
x"078583c1",
x"83c107c2",
x"fcf41d23",
x"fda45783",
x"471d8b9d",
x"0ae78663",
x"4863471d",
x"47190cf7",
x"0cf74563",
x"d8634715",
x"470906e7",
x"00f74563",
x"0007d963",
x"8713a85d",
x"4785ffd7",
x"0ae7e763",
x"1783a035",
x"878dfda4",
x"87c107c2",
x"83c107c2",
x"07378b8d",
x"07138000",
x"078a0247",
x"439c97ba",
x"fef42023",
x"24234791",
x"a049fef4",
x"fda41783",
x"07c2878d",
x"07c287c1",
x"8b8d83c1",
x"80000737",
x"03470713",
x"97ba078a",
x"2023439c",
x"47a1fef4",
x"fef42423",
x"1783a8a1",
x"878dfda4",
x"87c107c2",
x"83c107c2",
x"07378b8d",
x"07138000",
x"078a0447",
x"439c97ba",
x"fef42023",
x"242347a1",
x"a03dfef4",
x"fda41783",
x"07c2878d",
x"07c287c1",
x"8b8d83c1",
x"80000737",
x"05470713",
x"97ba078a",
x"2023439c",
x"47a1fef4",
x"fef42423",
x"0001a011",
x"fec42703",
x"fe842783",
x"078597ba",
x"fdc42703",
x"e8e7e9e3",
x"fdc42783",
x"2e230785",
x"a829fcf4",
x"fd442703",
x"fec42783",
x"802397ba",
x"27830007",
x"0785fec4",
x"fef42623",
x"fec42703",
x"fdc42783",
x"fef760e3",
x"00010001",
x"61455432",
x"71798082",
x"1800d622",
x"0fa387aa",
x"4783fcf4",
x"b793fdf4",
x"b7930307",
x"f7130017",
x"47830ff7",
x"b793fdf4",
x"f79303a7",
x"8ff90ff7",
x"0ff7f793",
x"fef407a3",
x"fef44783",
x"5432853e",
x"80826145",
x"d6067179",
x"1800d422",
x"fca42e23",
x"fcb42c23",
x"fdc42783",
x"2623439c",
x"2423fef4",
x"ac3dfe04",
x"fec42783",
x"0007c783",
x"fef403a3",
x"fe744703",
x"02c00793",
x"00f71863",
x"fec42783",
x"26230785",
x"a43dfef4",
x"fe842703",
x"ed63479d",
x"27831ee7",
x"9713fe84",
x"67a10027",
x"42478793",
x"439c97ba",
x"47838782",
x"853efe74",
x"87aa3fa9",
x"4791c789",
x"fef42423",
x"4703a0a1",
x"0793fe74",
x"086302b0",
x"470300f7",
x"0793fe74",
x"166302d0",
x"478900f7",
x"fef42423",
x"4703a025",
x"0793fe74",
x"166302e0",
x"479500f7",
x"fef42423",
x"4785a811",
x"fef42423",
x"fd842783",
x"43980791",
x"c3980705",
x"fd842783",
x"8713439c",
x"27830017",
x"c398fd84",
x"4783a259",
x"853efe74",
x"87aa35fd",
x"4791cb99",
x"fef42423",
x"fd842783",
x"439807a1",
x"c3980705",
x"4703a29d",
x"0793fe74",
x"1c6302e0",
x"479500f7",
x"fef42423",
x"fd842783",
x"439807a1",
x"c3980705",
x"4785a299",
x"fef42423",
x"fd842783",
x"439807a1",
x"c3980705",
x"4703aa0d",
x"0793fe74",
x"1c6302e0",
x"479500f7",
x"fef42423",
x"fd842783",
x"439807c1",
x"c3980705",
x"4783a221",
x"853efe74",
x"87aa3dad",
x"0e079e63",
x"24234785",
x"2783fef4",
x"07c1fd84",
x"07054398",
x"a0ddc398",
x"fe744703",
x"04500793",
x"00f70863",
x"fe744703",
x"06500793",
x"00f71c63",
x"2423478d",
x"2783fef4",
x"07d1fd84",
x"07054398",
x"a87dc398",
x"fe744783",
x"3535853e",
x"ebcd87aa",
x"24234785",
x"2783fef4",
x"07d1fd84",
x"07054398",
x"a879c398",
x"fe744703",
x"02b00793",
x"00f70863",
x"fe744703",
x"02d00793",
x"00f71c63",
x"24234799",
x"2783fef4",
x"07b1fd84",
x"07054398",
x"a8a5c398",
x"24234785",
x"2783fef4",
x"07b1fd84",
x"07054398",
x"a095c398",
x"fe744783",
x"33f1853e",
x"cb9987aa",
x"2423479d",
x"2783fef4",
x"07e1fd84",
x"07054398",
x"a091c398",
x"24234785",
x"2783fef4",
x"07e1fd84",
x"07054398",
x"a805c398",
x"fe744783",
x"3b61853e",
x"e38d87aa",
x"24234785",
x"2783fef4",
x"0791fd84",
x"07054398",
x"a039c398",
x"a0310001",
x"a0210001",
x"a0110001",
x"27830001",
x"0785fec4",
x"fef42623",
x"fec42783",
x"0007c783",
x"2703c791",
x"4785fe84",
x"daf71ae3",
x"fdc42783",
x"fec42703",
x"2783c398",
x"853efe84",
x"542250b2",
x"80826145",
x"d6227179",
x"2e231800",
x"2703fca4",
x"4795fdc4",
x"04e7eb63",
x"fdc42783",
x"00279713",
x"879367a1",
x"97ba4447",
x"8782439c",
x"800007b7",
x"0787a783",
x"fef42623",
x"a783a825",
x"26238141",
x"a03dfef4",
x"800007b7",
x"0687a783",
x"fef42623",
x"07b7a005",
x"a7838000",
x"262306c7",
x"a809fef4",
x"8181a783",
x"fef42623",
x"2623a021",
x"0001fe04",
x"fec42783",
x"5432853e",
x"80826145",
x"ce221101",
x"26231000",
x"2783fea4",
x"a073fec4",
x"00013007",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"3047a073",
x"44720001",
x"80826105",
x"ce061101",
x"1000cc22",
x"fea42623",
x"feb42423",
x"fec42783",
x"04278793",
x"fe842583",
x"38e1853e",
x"40f20001",
x"61054462",
x"11018082",
x"cc22ce06",
x"26231000",
x"2423fea4",
x"2783feb4",
x"8793fec4",
x"25830427",
x"853efe84",
x"000132a9",
x"446240f2",
x"80826105",
x"d6867159",
x"1880d4a2",
x"d0ef4509",
x"2423a5af",
x"d0effea4",
x"67f1a8af",
x"20078593",
x"fe842503",
x"fb4fd0ef",
x"e24fd0ef",
x"fe042623",
x"67ada829",
x"38a78593",
x"fec42503",
x"e4afd0ef",
x"fec42783",
x"26230785",
x"2703fef4",
x"47bdfec4",
x"fee7f1e3",
x"08018513",
x"862fe0ef",
x"859367ad",
x"451d3347",
x"dfcfd0ef",
x"b62fd0ef",
x"86ae862a",
x"05136531",
x"45813505",
x"00a60733",
x"3833883a",
x"87b300c8",
x"06b300b6",
x"87b600f8",
x"85be853a",
x"b16fd0ef",
x"08000513",
x"45213dfd",
x"67a535c5",
x"79278793",
x"fef42223",
x"f9c40793",
x"fe842583",
x"3dfd853e",
x"f9c40713",
x"fe442783",
x"fe842583",
x"9782853a",
x"fea42023",
x"f9c40793",
x"fe042583",
x"3721853e",
x"bfc90001",
x"ce221101",
x"27f31000",
x"26233000",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"341027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce221101",
x"27f31000",
x"26233430",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"34a027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"c6061141",
x"0800c422",
x"800007b7",
x"00078713",
x"87936785",
x"85bedea7",
x"c0ef853a",
x"d0efd3bf",
x"862aa2ef",
x"c53786ae",
x"05130578",
x"45811c05",
x"00a60733",
x"3833883a",
x"87b300c8",
x"06b300b6",
x"87b600f8",
x"85be853a",
x"a1efd0ef",
x"40b20001",
x"01414422",
x"71698082",
x"12112623",
x"12812423",
x"3f1d1a00",
x"fea42623",
x"fec42583",
x"08018513",
x"f7dfd0ef",
x"a64fd0ef",
x"fea42423",
x"fe842583",
x"08018513",
x"f69fd0ef",
x"fe842703",
x"800007b7",
x"ff6307bd",
x"270300e7",
x"07b7fe84",
x"07fd8000",
x"00e7e863",
x"85134585",
x"d0ef0801",
x"a039f43f",
x"0ff00593",
x"08018513",
x"f35fd0ef",
x"22233ddd",
x"2583fea4",
x"8513fe44",
x"d0ef0801",
x"3f21f23f",
x"fea42023",
x"fe042583",
x"08018513",
x"f11fd0ef",
x"2e2335f5",
x"2583fca4",
x"8513fdc4",
x"d0ef0801",
x"0713efff",
x"8613ed44",
x"45c10801",
x"d0ef853a",
x"0793d05f",
x"853eed44",
x"dc5fd0ef",
x"10500073",
x"0000bff5",
x"3340d4b0",
x"e7146a79",
x"0000e3c1",
x"1199be52",
x"1fd75608",
x"00000747",
x"39bf5e47",
x"8e3ae5a4",
x"00008d84",
x"00008374",
x"0000837c",
x"00008384",
x"0000838c",
x"00008394",
x"000083a0",
x"000083ac",
x"000083b8",
x"000083c4",
x"000083d0",
x"000083dc",
x"000083e8",
x"000083f4",
x"00008400",
x"0000840c",
x"00008418",
x"00000000",
x"00000066",
x"0000001e",
x"00000001"
);
end neorv32_application_image;

-- #################################################################################################
-- # << NEORV32 - Main VHDL Package File (CPU and SoC) >>                                          #
-- # ********************************************************************************************* #
-- # BSD 3-Clause License                                                                          #
-- #                                                                                               #
-- # Copyright (c) 2023, Stephan Nolting. All rights reserved.                                     #
-- #                                                                                               #
-- # Redistribution and use in source and binary forms, with or without modification, are          #
-- # permitted provided that the following conditions are met:                                     #
-- #                                                                                               #
-- # 1. Redistributions of source code must retain the above copyright notice, this list of        #
-- #    conditions and the following disclaimer.                                                   #
-- #                                                                                               #
-- # 2. Redistributions in binary form must reproduce the above copyright notice, this list of     #
-- #    conditions and the following disclaimer in the documentation and/or other materials        #
-- #    provided with the distribution.                                                            #
-- #                                                                                               #
-- # 3. Neither the name of the copyright holder nor the names of its contributors may be used to  #
-- #    endorse or promote products derived from this software without specific prior written      #
-- #    permission.                                                                                #
-- #                                                                                               #
-- # THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS   #
-- # OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF               #
-- # MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE    #
-- # COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL,     #
-- # EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE #
-- # GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED    #
-- # AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING     #
-- # NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED  #
-- # OF THE POSSIBILITY OF SUCH DAMAGE.                                                            #
-- # ********************************************************************************************* #
-- # The NEORV32 RISC-V Processor - https://github.com/stnolting/neorv32       (c) Stephan Nolting #
-- #################################################################################################

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package neorv32_package is

-- ****************************************************************************************************************************
-- Architecture Configuration and Constants
-- ****************************************************************************************************************************

  -- Architecture Configuration -------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- max response time for processor-internal bus transactions --
  -- = cycles after which an *unacknowledged* internal bus access will timeout triggering a bus fault exception
  constant bus_timeout_c : natural := 15; -- default = 15

  -- instruction prefetch buffer depth --
  constant ipb_depth_c : natural := 2; -- hast to be a power of two, min 2, default 2

  -- instruction monitor: raise exception if multi-cycle operation times out --
  constant monitor_mc_tmo_c : natural := 9; -- = log2 of max execution cycles (default = 512 cycles)

  -- Architecture Constants -----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant hw_version_c : std_ulogic_vector(31 downto 0) := x"01090200"; -- hardware version
  constant archid_c     : natural := 19; -- official RISC-V architecture ID
  constant XLEN         : natural := 32; -- native data path width, do not change!

  -- Check if we're inside the Matrix -------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant is_simulation_c : boolean := false -- seems like we're on real hardware
-- pragma translate_off
-- synthesis translate_off
-- RTL_SYNTHESIS OFF
  or true -- this MIGHT be a simulation
-- RTL_SYNTHESIS ON
-- synthesis translate_on
-- pragma translate_on
  ;

-- ****************************************************************************************************************************
-- Processor Address Space Layout
-- ****************************************************************************************************************************

  -- Main Address Regions ---
  constant mem_imem_base_c : std_ulogic_vector(31 downto 0) := x"00000000"; -- IMEM size via generic
  constant mem_dmem_base_c : std_ulogic_vector(31 downto 0) := x"80000000"; -- DMEM size via generic
  constant mem_xip_base_c  : std_ulogic_vector(31 downto 0) := x"e0000000"; -- page (4MSBs) only!
  constant mem_xip_size_c  : natural := 256*1024*1024;
  constant mem_boot_base_c : std_ulogic_vector(31 downto 0) := x"ffffc000";
  constant mem_boot_size_c : natural := 8*1024;
  constant mem_io_base_c   : std_ulogic_vector(31 downto 0) := x"ffffe000";
  constant mem_io_size_c   : natural := 8*1024;

  -- Start of uncached memory access (256MB page / 4MSBs only) --
  constant uncached_begin_c  : std_ulogic_vector(31 downto 0) := x"f0000000";

  -- IO Address Map --
  constant iodev_size_c      : natural := 256; -- size of a single IO device (bytes)
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe000"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe100"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe200"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe300"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe400"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe500"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe600"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe700"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe800"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffe900"; -- reserved
--constant base_io_???_c     : std_ulogic_vector(31 downto 0) := x"ffffea00"; -- reserved
  constant base_io_cfs_c     : std_ulogic_vector(31 downto 0) := x"ffffeb00";
  constant base_io_slink_c   : std_ulogic_vector(31 downto 0) := x"ffffec00";
  constant base_io_dma_c     : std_ulogic_vector(31 downto 0) := x"ffffed00";
  constant base_io_crc_c     : std_ulogic_vector(31 downto 0) := x"ffffee00";
  constant base_io_xip_c     : std_ulogic_vector(31 downto 0) := x"ffffef00";
  constant base_io_pwm_c     : std_ulogic_vector(31 downto 0) := x"fffff000";
  constant base_io_gptmr_c   : std_ulogic_vector(31 downto 0) := x"fffff100";
  constant base_io_onewire_c : std_ulogic_vector(31 downto 0) := x"fffff200";
  constant base_io_xirq_c    : std_ulogic_vector(31 downto 0) := x"fffff300";
  constant base_io_mtime_c   : std_ulogic_vector(31 downto 0) := x"fffff400";
  constant base_io_uart0_c   : std_ulogic_vector(31 downto 0) := x"fffff500";
  constant base_io_uart1_c   : std_ulogic_vector(31 downto 0) := x"fffff600";
  constant base_io_sdi_c     : std_ulogic_vector(31 downto 0) := x"fffff700";
  constant base_io_spi_c     : std_ulogic_vector(31 downto 0) := x"fffff800";
  constant base_io_twi_c     : std_ulogic_vector(31 downto 0) := x"fffff900";
  constant base_io_trng_c    : std_ulogic_vector(31 downto 0) := x"fffffa00";
  constant base_io_wdt_c     : std_ulogic_vector(31 downto 0) := x"fffffb00";
  constant base_io_gpio_c    : std_ulogic_vector(31 downto 0) := x"fffffc00";
  constant base_io_neoled_c  : std_ulogic_vector(31 downto 0) := x"fffffd00";
  constant base_io_sysinfo_c : std_ulogic_vector(31 downto 0) := x"fffffe00";
  constant base_io_dm_c      : std_ulogic_vector(31 downto 0) := x"ffffff00";

  -- On-Chip Debugger - Debug Module Entry Points (Code ROM) --
  constant dm_exc_entry_c  : std_ulogic_vector(31 downto 0) := x"ffffff00"; -- = base_io_dm_c + 0, exceptions entry point
  constant dm_park_entry_c : std_ulogic_vector(31 downto 0) := x"ffffff08"; -- = base_io_dm_c + 8, normal entry point

-- ****************************************************************************************************************************
-- SoC Definitions
-- ****************************************************************************************************************************

  -- SoC Clock Select -----------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant clk_div2_c    : natural := 0;
  constant clk_div4_c    : natural := 1;
  constant clk_div8_c    : natural := 2;
  constant clk_div64_c   : natural := 3;
  constant clk_div128_c  : natural := 4;
  constant clk_div1024_c : natural := 5;
  constant clk_div2048_c : natural := 6;
  constant clk_div4096_c : natural := 7;

  -- Internal Memory Types ------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  type mem32_t is array (natural range <>) of std_ulogic_vector(31 downto 0); -- memory with 32-bit entries
  type mem16_t is array (natural range <>) of std_ulogic_vector(15 downto 0); -- memory with 16-bit entries
  type mem8_t  is array (natural range <>) of std_ulogic_vector(07 downto 0); -- memory with 8-bit entries
  
  type mem15_t  is array (natural range <>) of std_ulogic_vector(14 downto 0); -- memory with 15-bit entries
  type mem13_t  is array (natural range <>) of std_ulogic_vector(12 downto 0); -- memory with 13-bit entries

  -- Internal Bus Interface -----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- bus request --
  type bus_req_t is record
    addr : std_ulogic_vector(31 downto 0); -- access address
    data : std_ulogic_vector(31 downto 0); -- write data
    ben  : std_ulogic_vector(03 downto 0); -- byte enable
    stb  : std_ulogic; -- request strobe (single-shot)
    rw   : std_ulogic; -- 0=read, 1=write
    src  : std_ulogic; -- access source (1=instruction fetch, 0=data access)
    priv : std_ulogic; -- set if privileged (machine-mode) access
    rvso : std_ulogic; -- set if reservation set operation (atomic LR/SC)
  end record;

  -- bus response --
  type bus_rsp_t is record
    data : std_ulogic_vector(31 downto 0); -- read data
    ack  : std_ulogic; -- access acknowledge (single-shot)
    err  : std_ulogic; -- access error (single-shot)
  end record;

  -- source (request) termination --
  constant req_terminate_c : bus_req_t := (
    addr => (others => '0'),
    data => (others => '0'),
    ben  => (others => '0'),
    stb  => '0',
    rw   => '0',
    src  => '0',
    priv => '0',
    rvso => '0'
  );

  -- endpoint (response) termination --
  constant rsp_terminate_c : bus_rsp_t := (
    data => (others => '0'),
    ack  => '0',
    err  => '0'
  );

  -- Debug Module Interface -----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- request --
  type dmi_req_t is record
    addr : std_ulogic_vector(06 downto 0);
    op   : std_ulogic_vector(01 downto 0);
    data : std_ulogic_vector(31 downto 0);
  end record;

  -- request operation --
  constant dmi_req_nop_c : std_ulogic_vector(1 downto 0) := "00"; -- no operation
  constant dmi_req_rd_c  : std_ulogic_vector(1 downto 0) := "01"; -- read access
  constant dmi_req_wr_c  : std_ulogic_vector(1 downto 0) := "10"; -- write access

  -- response --
  type dmi_rsp_t is record
    data : std_ulogic_vector(31 downto 0);
    ack  : std_ulogic;
  end record;

-- ****************************************************************************************************************************
-- RISC-V ISA Definitions
-- ****************************************************************************************************************************

  -- RISC-V 32-Bit Instruction Word Layout --------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant instr_opcode_lsb_c  : natural :=  0; -- opcode bit 0
  constant instr_opcode_msb_c  : natural :=  6; -- opcode bit 6
  constant instr_rd_lsb_c      : natural :=  7; -- destination register address bit 0
  constant instr_rd_msb_c      : natural := 11; -- destination register address bit 4
  constant instr_funct3_lsb_c  : natural := 12; -- funct3 bit 0
  constant instr_funct3_msb_c  : natural := 14; -- funct3 bit 2
  constant instr_rs1_lsb_c     : natural := 15; -- source register 1 address bit 0
  constant instr_rs1_msb_c     : natural := 19; -- source register 1 address bit 4
  constant instr_rs2_lsb_c     : natural := 20; -- source register 2 address bit 0
  constant instr_rs2_msb_c     : natural := 24; -- source register 2 address bit 4
  constant instr_rs3_lsb_c     : natural := 27; -- source register 3 address bit 0
  constant instr_rs3_msb_c     : natural := 31; -- source register 3 address bit 4
  constant instr_funct7_lsb_c  : natural := 25; -- funct7 bit 0
  constant instr_funct7_msb_c  : natural := 31; -- funct7 bit 6
  constant instr_funct12_lsb_c : natural := 20; -- funct12 bit 0
  constant instr_funct12_msb_c : natural := 31; -- funct12 bit 11
  constant instr_imm12_lsb_c   : natural := 20; -- immediate12 bit 0
  constant instr_imm12_msb_c   : natural := 31; -- immediate12 bit 11
  constant instr_imm20_lsb_c   : natural := 12; -- immediate20 bit 0
  constant instr_imm20_msb_c   : natural := 31; -- immediate20 bit 21
  constant instr_funct5_lsb_c  : natural := 27; -- funct5 select bit 0
  constant instr_funct5_msb_c  : natural := 31; -- funct5 select bit 4

  -- RISC-V Opcodes -------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- alu --
  constant opcode_alui_c   : std_ulogic_vector(6 downto 0) := "0010011"; -- ALU operation with immediate
  constant opcode_alu_c    : std_ulogic_vector(6 downto 0) := "0110011"; -- ALU operation
  constant opcode_lui_c    : std_ulogic_vector(6 downto 0) := "0110111"; -- load upper immediate
  constant opcode_auipc_c  : std_ulogic_vector(6 downto 0) := "0010111"; -- add upper immediate to PC
  -- control flow --
  constant opcode_jal_c    : std_ulogic_vector(6 downto 0) := "1101111"; -- jump and link
  constant opcode_jalr_c   : std_ulogic_vector(6 downto 0) := "1100111"; -- jump and link with register
  constant opcode_branch_c : std_ulogic_vector(6 downto 0) := "1100011"; -- branch
  -- memory access --
  constant opcode_load_c   : std_ulogic_vector(6 downto 0) := "0000011"; -- load
  constant opcode_store_c  : std_ulogic_vector(6 downto 0) := "0100011"; -- store
  constant opcode_amo_c    : std_ulogic_vector(6 downto 0) := "0101111"; -- atomic memory access
  constant opcode_fence_c  : std_ulogic_vector(6 downto 0) := "0001111"; -- fence / fence.i
  -- system/csr --
  constant opcode_system_c : std_ulogic_vector(6 downto 0) := "1110011"; -- system/csr access
  -- floating point operations --
  constant opcode_fop_c    : std_ulogic_vector(6 downto 0) := "1010011"; -- dual/single operand instruction
  -- official custom RISC-V opcodes - free for custom instructions --
  constant opcode_cust0_c  : std_ulogic_vector(6 downto 0) := "0001011"; -- custom-0
  constant opcode_cust1_c  : std_ulogic_vector(6 downto 0) := "0101011"; -- custom-1
  constant opcode_cust2_c  : std_ulogic_vector(6 downto 0) := "1011011"; -- custom-2
  constant opcode_cust3_c  : std_ulogic_vector(6 downto 0) := "1111011"; -- custom-3

  -- RISC-V Funct3 --------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- control flow --
  constant funct3_beq_c    : std_ulogic_vector(2 downto 0) := "000"; -- branch if equal
  constant funct3_bne_c    : std_ulogic_vector(2 downto 0) := "001"; -- branch if not equal
  constant funct3_blt_c    : std_ulogic_vector(2 downto 0) := "100"; -- branch if less than
  constant funct3_bge_c    : std_ulogic_vector(2 downto 0) := "101"; -- branch if greater than or equal
  constant funct3_bltu_c   : std_ulogic_vector(2 downto 0) := "110"; -- branch if less than (unsigned)
  constant funct3_bgeu_c   : std_ulogic_vector(2 downto 0) := "111"; -- branch if greater than or equal (unsigned)
  -- memory access --
  constant funct3_lb_c     : std_ulogic_vector(2 downto 0) := "000"; -- load byte (signed)
  constant funct3_lh_c     : std_ulogic_vector(2 downto 0) := "001"; -- load half word (signed)
  constant funct3_lw_c     : std_ulogic_vector(2 downto 0) := "010"; -- load word (signed)
  constant funct3_lbu_c    : std_ulogic_vector(2 downto 0) := "100"; -- load byte (unsigned)
  constant funct3_lhu_c    : std_ulogic_vector(2 downto 0) := "101"; -- load half word (unsigned)
  constant funct3_lwu_c    : std_ulogic_vector(2 downto 0) := "110"; -- load word (unsigned)
  constant funct3_sb_c     : std_ulogic_vector(2 downto 0) := "000"; -- store byte
  constant funct3_sh_c     : std_ulogic_vector(2 downto 0) := "001"; -- store half word
  constant funct3_sw_c     : std_ulogic_vector(2 downto 0) := "010"; -- store word
  -- alu --
  constant funct3_subadd_c : std_ulogic_vector(2 downto 0) := "000"; -- sub/add via funct7
  constant funct3_sll_c    : std_ulogic_vector(2 downto 0) := "001"; -- shift logical left
  constant funct3_slt_c    : std_ulogic_vector(2 downto 0) := "010"; -- set on less
  constant funct3_sltu_c   : std_ulogic_vector(2 downto 0) := "011"; -- set on less unsigned
  constant funct3_xor_c    : std_ulogic_vector(2 downto 0) := "100"; -- xor
  constant funct3_sr_c     : std_ulogic_vector(2 downto 0) := "101"; -- shift right via funct7
  constant funct3_or_c     : std_ulogic_vector(2 downto 0) := "110"; -- or
  constant funct3_and_c    : std_ulogic_vector(2 downto 0) := "111"; -- and
  -- system/csr --
  constant funct3_env_c    : std_ulogic_vector(2 downto 0) := "000"; -- ecall, ebreak, mret, wfi, ...
  constant funct3_csrrw_c  : std_ulogic_vector(2 downto 0) := "001"; -- csr r/w
  constant funct3_csrrs_c  : std_ulogic_vector(2 downto 0) := "010"; -- csr read & set
  constant funct3_csrrc_c  : std_ulogic_vector(2 downto 0) := "011"; -- csr read & clear
  constant funct3_csril_c  : std_ulogic_vector(2 downto 0) := "100"; -- undefined/illegal csr command
  constant funct3_csrrwi_c : std_ulogic_vector(2 downto 0) := "101"; -- csr r/w immediate
  constant funct3_csrrsi_c : std_ulogic_vector(2 downto 0) := "110"; -- csr read & set immediate
  constant funct3_csrrci_c : std_ulogic_vector(2 downto 0) := "111"; -- csr read & clear immediate
  -- fence --
  constant funct3_fence_c  : std_ulogic_vector(2 downto 0) := "000"; -- fence - order IO/memory access
  constant funct3_fencei_c : std_ulogic_vector(2 downto 0) := "001"; -- fence.i - instruction stream sync

  -- RISC-V Funct12 - SYSTEM ----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant funct12_ecall_c  : std_ulogic_vector(11 downto 0) := x"000"; -- ecall
  constant funct12_ebreak_c : std_ulogic_vector(11 downto 0) := x"001"; -- ebreak
  constant funct12_wfi_c    : std_ulogic_vector(11 downto 0) := x"105"; -- wfi
  constant funct12_mret_c   : std_ulogic_vector(11 downto 0) := x"302"; -- mret
  constant funct12_dret_c   : std_ulogic_vector(11 downto 0) := x"7b2"; -- dret

  -- RISC-V Floating-Point Stuff ------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant float_single_c : std_ulogic_vector(1 downto 0) := "00"; -- single-precision (32-bit)
--constant float_double_c : std_ulogic_vector(1 downto 0) := "01"; -- double-precision (64-bit)
--constant float_half_c   : std_ulogic_vector(1 downto 0) := "10"; -- half-precision (16-bit)
--constant float_quad_c   : std_ulogic_vector(1 downto 0) := "11"; -- quad-precision (128-bit)

  -- number class flags --
  constant fp_class_neg_inf_c    : natural := 0; -- negative infinity
  constant fp_class_neg_norm_c   : natural := 1; -- negative normal number
  constant fp_class_neg_denorm_c : natural := 2; -- negative subnormal number
  constant fp_class_neg_zero_c   : natural := 3; -- negative zero
  constant fp_class_pos_zero_c   : natural := 4; -- positive zero
  constant fp_class_pos_denorm_c : natural := 5; -- positive subnormal number
  constant fp_class_pos_norm_c   : natural := 6; -- positive normal number
  constant fp_class_pos_inf_c    : natural := 7; -- positive infinity
  constant fp_class_snan_c       : natural := 8; -- signaling NaN (sNaN)
  constant fp_class_qnan_c       : natural := 9; -- quiet NaN (qNaN)

  -- exception flags --
  constant fp_exc_nx_c : natural := 0; -- inexact
  constant fp_exc_uf_c : natural := 1; -- underflow
  constant fp_exc_of_c : natural := 2; -- overflow
  constant fp_exc_dz_c : natural := 3; -- division by zero
  constant fp_exc_nv_c : natural := 4; -- invalid operation

  -- special values (single-precision) --
  constant fp_single_qnan_c     : std_ulogic_vector(31 downto 0) := x"7fc00000"; -- quiet NaN
  constant fp_single_snan_c     : std_ulogic_vector(31 downto 0) := x"7fa00000"; -- signaling NaN
  constant fp_single_pos_inf_c  : std_ulogic_vector(31 downto 0) := x"7f800000"; -- positive infinity
  constant fp_single_neg_inf_c  : std_ulogic_vector(31 downto 0) := x"ff800000"; -- negative infinity
  constant fp_single_pos_zero_c : std_ulogic_vector(31 downto 0) := x"00000000"; -- positive zero
  constant fp_single_neg_zero_c : std_ulogic_vector(31 downto 0) := x"80000000"; -- negative zero

  -- RISC-V CSRs ----------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- user floating-point CSRs --
  constant csr_fflags_c         : std_ulogic_vector(11 downto 0) := x"001";
  constant csr_frm_c            : std_ulogic_vector(11 downto 0) := x"002";
  constant csr_fcsr_c           : std_ulogic_vector(11 downto 0) := x"003";
  -- machine trap setup --
  constant csr_mstatus_c        : std_ulogic_vector(11 downto 0) := x"300";
  constant csr_misa_c           : std_ulogic_vector(11 downto 0) := x"301";
  constant csr_mie_c            : std_ulogic_vector(11 downto 0) := x"304";
  constant csr_mtvec_c          : std_ulogic_vector(11 downto 0) := x"305";
  constant csr_mcounteren_c     : std_ulogic_vector(11 downto 0) := x"306";
  constant csr_mstatush_c       : std_ulogic_vector(11 downto 0) := x"310";
  -- machine configuration --
  constant csr_menvcfg_c        : std_ulogic_vector(11 downto 0) := x"30a";
  constant csr_menvcfgh_c       : std_ulogic_vector(11 downto 0) := x"31a";
  -- machine counter setup --
  constant csr_mcountinhibit_c  : std_ulogic_vector(11 downto 0) := x"320";
  constant csr_mcyclecfg_c      : std_ulogic_vector(11 downto 0) := x"321";
  constant csr_minstretcfg_c    : std_ulogic_vector(11 downto 0) := x"322";
  constant csr_mhpmevent3_c     : std_ulogic_vector(11 downto 0) := x"323";
  constant csr_mhpmevent4_c     : std_ulogic_vector(11 downto 0) := x"324";
  constant csr_mhpmevent5_c     : std_ulogic_vector(11 downto 0) := x"325";
  constant csr_mhpmevent6_c     : std_ulogic_vector(11 downto 0) := x"326";
  constant csr_mhpmevent7_c     : std_ulogic_vector(11 downto 0) := x"327";
  constant csr_mhpmevent8_c     : std_ulogic_vector(11 downto 0) := x"328";
  constant csr_mhpmevent9_c     : std_ulogic_vector(11 downto 0) := x"329";
  constant csr_mhpmevent10_c    : std_ulogic_vector(11 downto 0) := x"32a";
  constant csr_mhpmevent11_c    : std_ulogic_vector(11 downto 0) := x"32b";
  constant csr_mhpmevent12_c    : std_ulogic_vector(11 downto 0) := x"32c";
  constant csr_mhpmevent13_c    : std_ulogic_vector(11 downto 0) := x"32d";
  constant csr_mhpmevent14_c    : std_ulogic_vector(11 downto 0) := x"32e";
  constant csr_mhpmevent15_c    : std_ulogic_vector(11 downto 0) := x"32f";
  -- machine trap handling --
  constant csr_mscratch_c       : std_ulogic_vector(11 downto 0) := x"340";
  constant csr_mepc_c           : std_ulogic_vector(11 downto 0) := x"341";
  constant csr_mcause_c         : std_ulogic_vector(11 downto 0) := x"342";
  constant csr_mtval_c          : std_ulogic_vector(11 downto 0) := x"343";
  constant csr_mip_c            : std_ulogic_vector(11 downto 0) := x"344";
  constant csr_mtinst_c         : std_ulogic_vector(11 downto 0) := x"34a";
  -- physical memory protection - configuration --
  constant csr_pmpcfg0_c        : std_ulogic_vector(11 downto 0) := x"3a0";
  constant csr_pmpcfg1_c        : std_ulogic_vector(11 downto 0) := x"3a1";
  constant csr_pmpcfg2_c        : std_ulogic_vector(11 downto 0) := x"3a2";
  constant csr_pmpcfg3_c        : std_ulogic_vector(11 downto 0) := x"3a3";
  -- physical memory protection - address --
  constant csr_pmpaddr0_c       : std_ulogic_vector(11 downto 0) := x"3b0";
  constant csr_pmpaddr1_c       : std_ulogic_vector(11 downto 0) := x"3b1";
  constant csr_pmpaddr2_c       : std_ulogic_vector(11 downto 0) := x"3b2";
  constant csr_pmpaddr3_c       : std_ulogic_vector(11 downto 0) := x"3b3";
  constant csr_pmpaddr4_c       : std_ulogic_vector(11 downto 0) := x"3b4";
  constant csr_pmpaddr5_c       : std_ulogic_vector(11 downto 0) := x"3b5";
  constant csr_pmpaddr6_c       : std_ulogic_vector(11 downto 0) := x"3b6";
  constant csr_pmpaddr7_c       : std_ulogic_vector(11 downto 0) := x"3b7";
  constant csr_pmpaddr8_c       : std_ulogic_vector(11 downto 0) := x"3b8";
  constant csr_pmpaddr9_c       : std_ulogic_vector(11 downto 0) := x"3b9";
  constant csr_pmpaddr10_c      : std_ulogic_vector(11 downto 0) := x"3ba";
  constant csr_pmpaddr11_c      : std_ulogic_vector(11 downto 0) := x"3bb";
  constant csr_pmpaddr12_c      : std_ulogic_vector(11 downto 0) := x"3bc";
  constant csr_pmpaddr13_c      : std_ulogic_vector(11 downto 0) := x"3bd";
  constant csr_pmpaddr14_c      : std_ulogic_vector(11 downto 0) := x"3be";
  constant csr_pmpaddr15_c      : std_ulogic_vector(11 downto 0) := x"3bf";
  -- machine counter setup - continued --
  constant csr_mcyclecfgh_c     : std_ulogic_vector(11 downto 0) := x"721";
  constant csr_minstretcfgh_c   : std_ulogic_vector(11 downto 0) := x"722";
  -- trigger module registers --
  constant csr_tselect_c        : std_ulogic_vector(11 downto 0) := x"7a0";
  constant csr_tdata1_c         : std_ulogic_vector(11 downto 0) := x"7a1";
  constant csr_tdata2_c         : std_ulogic_vector(11 downto 0) := x"7a2";
  constant csr_tinfo_c          : std_ulogic_vector(11 downto 0) := x"7a4";
  -- debug mode registers --
  constant csr_dcsr_c           : std_ulogic_vector(11 downto 0) := x"7b0";
  constant csr_dpc_c            : std_ulogic_vector(11 downto 0) := x"7b1";
  constant csr_dscratch0_c      : std_ulogic_vector(11 downto 0) := x"7b2";
  -- NEORV32-specific (user-mode) registers --
  constant csr_cfureg0_c        : std_ulogic_vector(11 downto 0) := x"800";
  constant csr_cfureg1_c        : std_ulogic_vector(11 downto 0) := x"801";
  constant csr_cfureg2_c        : std_ulogic_vector(11 downto 0) := x"802";
  constant csr_cfureg3_c        : std_ulogic_vector(11 downto 0) := x"803";
  -- machine counters/timers --
  constant csr_mcycle_c         : std_ulogic_vector(11 downto 0) := x"b00";
--constant csr_mtime_c          : std_ulogic_vector(11 downto 0) := x"b01";
  constant csr_minstret_c       : std_ulogic_vector(11 downto 0) := x"b02";
  constant csr_mhpmcounter3_c   : std_ulogic_vector(11 downto 0) := x"b03";
  constant csr_mhpmcounter4_c   : std_ulogic_vector(11 downto 0) := x"b04";
  constant csr_mhpmcounter5_c   : std_ulogic_vector(11 downto 0) := x"b05";
  constant csr_mhpmcounter6_c   : std_ulogic_vector(11 downto 0) := x"b06";
  constant csr_mhpmcounter7_c   : std_ulogic_vector(11 downto 0) := x"b07";
  constant csr_mhpmcounter8_c   : std_ulogic_vector(11 downto 0) := x"b08";
  constant csr_mhpmcounter9_c   : std_ulogic_vector(11 downto 0) := x"b09";
  constant csr_mhpmcounter10_c  : std_ulogic_vector(11 downto 0) := x"b0a";
  constant csr_mhpmcounter11_c  : std_ulogic_vector(11 downto 0) := x"b0b";
  constant csr_mhpmcounter12_c  : std_ulogic_vector(11 downto 0) := x"b0c";
  constant csr_mhpmcounter13_c  : std_ulogic_vector(11 downto 0) := x"b0d";
  constant csr_mhpmcounter14_c  : std_ulogic_vector(11 downto 0) := x"b0e";
  constant csr_mhpmcounter15_c  : std_ulogic_vector(11 downto 0) := x"b0f";
  --
  constant csr_mcycleh_c        : std_ulogic_vector(11 downto 0) := x"b80";
--constant csr_mtimeh_c         : std_ulogic_vector(11 downto 0) := x"b81";
  constant csr_minstreth_c      : std_ulogic_vector(11 downto 0) := x"b82";
  constant csr_mhpmcounter3h_c  : std_ulogic_vector(11 downto 0) := x"b83";
  constant csr_mhpmcounter4h_c  : std_ulogic_vector(11 downto 0) := x"b84";
  constant csr_mhpmcounter5h_c  : std_ulogic_vector(11 downto 0) := x"b85";
  constant csr_mhpmcounter6h_c  : std_ulogic_vector(11 downto 0) := x"b86";
  constant csr_mhpmcounter7h_c  : std_ulogic_vector(11 downto 0) := x"b87";
  constant csr_mhpmcounter8h_c  : std_ulogic_vector(11 downto 0) := x"b88";
  constant csr_mhpmcounter9h_c  : std_ulogic_vector(11 downto 0) := x"b89";
  constant csr_mhpmcounter10h_c : std_ulogic_vector(11 downto 0) := x"b8a";
  constant csr_mhpmcounter11h_c : std_ulogic_vector(11 downto 0) := x"b8b";
  constant csr_mhpmcounter12h_c : std_ulogic_vector(11 downto 0) := x"b8c";
  constant csr_mhpmcounter13h_c : std_ulogic_vector(11 downto 0) := x"b8d";
  constant csr_mhpmcounter14h_c : std_ulogic_vector(11 downto 0) := x"b8e";
  constant csr_mhpmcounter15h_c : std_ulogic_vector(11 downto 0) := x"b8f";
  -- user counters/timers --
  constant csr_cycle_c          : std_ulogic_vector(11 downto 0) := x"c00";
  constant csr_time_c           : std_ulogic_vector(11 downto 0) := x"c01";
  constant csr_instret_c        : std_ulogic_vector(11 downto 0) := x"c02";
  constant csr_hpmcounter3_c    : std_ulogic_vector(11 downto 0) := x"c03";
  constant csr_hpmcounter4_c    : std_ulogic_vector(11 downto 0) := x"c04";
  constant csr_hpmcounter5_c    : std_ulogic_vector(11 downto 0) := x"c05";
  constant csr_hpmcounter6_c    : std_ulogic_vector(11 downto 0) := x"c06";
  constant csr_hpmcounter7_c    : std_ulogic_vector(11 downto 0) := x"c07";
  constant csr_hpmcounter8_c    : std_ulogic_vector(11 downto 0) := x"c08";
  constant csr_hpmcounter9_c    : std_ulogic_vector(11 downto 0) := x"c09";
  constant csr_hpmcounter10_c   : std_ulogic_vector(11 downto 0) := x"c0a";
  constant csr_hpmcounter11_c   : std_ulogic_vector(11 downto 0) := x"c0b";
  constant csr_hpmcounter12_c   : std_ulogic_vector(11 downto 0) := x"c0c";
  constant csr_hpmcounter13_c   : std_ulogic_vector(11 downto 0) := x"c0d";
  constant csr_hpmcounter14_c   : std_ulogic_vector(11 downto 0) := x"c0e";
  constant csr_hpmcounter15_c   : std_ulogic_vector(11 downto 0) := x"c0f";
  --
  constant csr_cycleh_c         : std_ulogic_vector(11 downto 0) := x"c80";
  constant csr_timeh_c          : std_ulogic_vector(11 downto 0) := x"c81";
  constant csr_instreth_c       : std_ulogic_vector(11 downto 0) := x"c82";
  constant csr_hpmcounter3h_c   : std_ulogic_vector(11 downto 0) := x"c83";
  constant csr_hpmcounter4h_c   : std_ulogic_vector(11 downto 0) := x"c84";
  constant csr_hpmcounter5h_c   : std_ulogic_vector(11 downto 0) := x"c85";
  constant csr_hpmcounter6h_c   : std_ulogic_vector(11 downto 0) := x"c86";
  constant csr_hpmcounter7h_c   : std_ulogic_vector(11 downto 0) := x"c87";
  constant csr_hpmcounter8h_c   : std_ulogic_vector(11 downto 0) := x"c88";
  constant csr_hpmcounter9h_c   : std_ulogic_vector(11 downto 0) := x"c89";
  constant csr_hpmcounter10h_c  : std_ulogic_vector(11 downto 0) := x"c8a";
  constant csr_hpmcounter11h_c  : std_ulogic_vector(11 downto 0) := x"c8b";
  constant csr_hpmcounter12h_c  : std_ulogic_vector(11 downto 0) := x"c8c";
  constant csr_hpmcounter13h_c  : std_ulogic_vector(11 downto 0) := x"c8d";
  constant csr_hpmcounter14h_c  : std_ulogic_vector(11 downto 0) := x"c8e";
  constant csr_hpmcounter15h_c  : std_ulogic_vector(11 downto 0) := x"c8f";
  -- machine information registers --
  constant csr_mvendorid_c      : std_ulogic_vector(11 downto 0) := x"f11";
  constant csr_marchid_c        : std_ulogic_vector(11 downto 0) := x"f12";
  constant csr_mimpid_c         : std_ulogic_vector(11 downto 0) := x"f13";
  constant csr_mhartid_c        : std_ulogic_vector(11 downto 0) := x"f14";
  constant csr_mconfigptr_c     : std_ulogic_vector(11 downto 0) := x"f15";
  -- NEORV32-specific (machine-mode) registers --
  constant csr_mxisa_c          : std_ulogic_vector(11 downto 0) := x"fc0";

-- ****************************************************************************************************************************
-- CPU Control
-- ****************************************************************************************************************************

  -- Main CPU Control Bus -------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  type ctrl_bus_t is record
    -- register file --
    rf_wb_en     : std_ulogic; -- write back enable
    rf_rs1       : std_ulogic_vector(04 downto 0); -- source register 1 address
    rf_rs2       : std_ulogic_vector(04 downto 0); -- source register 2 address
    rf_rs3       : std_ulogic_vector(04 downto 0); -- source register 3 address
    rf_rd        : std_ulogic_vector(04 downto 0); -- destination register address
    rf_mux       : std_ulogic_vector(01 downto 0); -- input source select
    rf_zero_we   : std_ulogic;                     -- allow/force write access to x0
    -- alu --
    alu_op       : std_ulogic_vector(02 downto 0); -- ALU operation select
    alu_opa_mux  : std_ulogic;                     -- operand A select (0=rs1, 1=PC)
    alu_opb_mux  : std_ulogic;                     -- operand B select (0=rs2, 1=IMM)
    alu_unsigned : std_ulogic;                     -- is unsigned ALU operation
    alu_cp_trig  : std_ulogic_vector(04 downto 0); -- co-processor trigger (one-hot)
    -- load/store unit --
    lsu_req      : std_ulogic;                     -- trigger memory access request
    lsu_rw       : std_ulogic;                     -- 0: read access, 1: write access
    lsu_mo_we    : std_ulogic;                     -- memory address and data output register write enable
    lsu_fence    : std_ulogic;                     -- fence operation
    lsu_fencei   : std_ulogic;                     -- fence.i operation
    lsu_priv     : std_ulogic;                     -- effective privilege level for load/store
    -- instruction word --
    ir_funct3    : std_ulogic_vector(02 downto 0); -- funct3 bit field
    ir_funct12   : std_ulogic_vector(11 downto 0); -- funct12 bit field
    ir_opcode    : std_ulogic_vector(06 downto 0); -- opcode bit field
    -- cpu status --
    cpu_priv     : std_ulogic;                     -- effective privilege mode
    cpu_sleep    : std_ulogic;                     -- set when CPU is in sleep mode
    cpu_trap     : std_ulogic;                     -- set when CPU is entering trap exec
    cpu_debug    : std_ulogic;                     -- set when CPU is in debug mode
  end record;

  -- control bus reset initializer --
  constant ctrl_bus_zero_c : ctrl_bus_t := (
    rf_wb_en     => '0',
    rf_rs1       => (others => '0'),
    rf_rs2       => (others => '0'),
    rf_rs3       => (others => '0'),
    rf_rd        => (others => '0'),
    rf_mux       => (others => '0'),
    rf_zero_we   => '0',
    alu_op       => (others => '0'),
    alu_opa_mux  => '0',
    alu_opb_mux  => '0',
    alu_unsigned => '0',
    alu_cp_trig  => (others => '0'),
    lsu_req      => '0',
    lsu_rw       => '0',
    lsu_mo_we    => '0',
    lsu_fence    => '0',
    lsu_fencei   => '0',
    lsu_priv     => '0',
    ir_funct3    => (others => '0'),
    ir_funct12   => (others => '0'),
    ir_opcode    => (others => '0'),
    cpu_priv     => '0',
    cpu_sleep    => '0',
    cpu_trap     => '0',
    cpu_debug    => '0'
  );

  -- Comparator Bus -------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant cmp_equal_c : natural := 0;
  constant cmp_less_c  : natural := 1; -- for signed and unsigned comparisons

  -- CPU Co-Processor IDs -------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant cp_sel_shifter_c  : natural := 0; -- CP0: shift operations (base ISA)
  constant cp_sel_muldiv_c   : natural := 1; -- CP1: multiplication/division operations ('M' extensions)
  constant cp_sel_bitmanip_c : natural := 2; -- CP2: bit manipulation ('B' extensions)
  constant cp_sel_fpu_c      : natural := 3; -- CP3: floating-point unit ('Zfinx' extension)
  constant cp_sel_cfu_c      : natural := 4; -- CP4: custom instructions CFU ('Zxcfu' extension)

  -- ALU Function Codes [DO NOT CHANGE ENCODING!] -------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant alu_op_add_c  : std_ulogic_vector(2 downto 0) := "000"; -- result <= A + B
  constant alu_op_sub_c  : std_ulogic_vector(2 downto 0) := "001"; -- result <= A - B
  constant alu_op_cp_c   : std_ulogic_vector(2 downto 0) := "010"; -- result <= ALU co-processor
  constant alu_op_slt_c  : std_ulogic_vector(2 downto 0) := "011"; -- result <= A < B
  constant alu_op_movb_c : std_ulogic_vector(2 downto 0) := "100"; -- result <= B
  constant alu_op_xor_c  : std_ulogic_vector(2 downto 0) := "101"; -- result <= A xor B
  constant alu_op_or_c   : std_ulogic_vector(2 downto 0) := "110"; -- result <= A or B
  constant alu_op_and_c  : std_ulogic_vector(2 downto 0) := "111"; -- result <= A and B

  -- Register File Input Select -------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant rf_mux_alu_c : std_ulogic_vector(1 downto 0) := "00"; -- register file <= alu result
  constant rf_mux_mem_c : std_ulogic_vector(1 downto 0) := "01"; -- register file <= memory read data
  constant rf_mux_csr_c : std_ulogic_vector(1 downto 0) := "10"; -- register file <= CSR read data
  constant rf_mux_ret_c : std_ulogic_vector(1 downto 0) := "11"; -- register file <= link-PC (return address)

  -- Trap ID Codes --------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- MSB:   1 = interrupt, 0 = sync. exception
  -- MSB-1: 1 = entry to debug mode, 0 = normal trapping
  -- RISC-V compliant synchronous exceptions --
  constant trap_ima_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00000"; -- 0: instruction misaligned
  constant trap_iaf_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00001"; -- 1: instruction access fault
  constant trap_iil_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00010"; -- 2: illegal instruction
  constant trap_brk_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00011"; -- 3: breakpoint
  constant trap_lma_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00100"; -- 4: load address misaligned
  constant trap_laf_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00101"; -- 5: load access fault
  constant trap_sma_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00110"; -- 6: store address misaligned
  constant trap_saf_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "00111"; -- 7: store access fault
  constant trap_env_c      : std_ulogic_vector(6 downto 0) := "0" & "0" & "010UU"; -- 8..11: environment call from u/s/h/m
  -- RISC-V compliant asynchronous exceptions (interrupts) --
  constant trap_msi_c      : std_ulogic_vector(6 downto 0) := "1" & "0" & "00011"; -- 3:  machine software interrupt
  constant trap_mti_c      : std_ulogic_vector(6 downto 0) := "1" & "0" & "00111"; -- 7:  machine timer interrupt
  constant trap_mei_c      : std_ulogic_vector(6 downto 0) := "1" & "0" & "01011"; -- 11: machine external interrupt
  -- NEORV32-specific (RISC-V custom) asynchronous exceptions (interrupts) --
  constant trap_firq0_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10000"; -- 16: fast interrupt 0
  constant trap_firq1_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10001"; -- 17: fast interrupt 1
  constant trap_firq2_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10010"; -- 18: fast interrupt 2
  constant trap_firq3_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10011"; -- 19: fast interrupt 3
  constant trap_firq4_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10100"; -- 20: fast interrupt 4
  constant trap_firq5_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10101"; -- 21: fast interrupt 5
  constant trap_firq6_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10110"; -- 22: fast interrupt 6
  constant trap_firq7_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "10111"; -- 23: fast interrupt 7
  constant trap_firq8_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "11000"; -- 24: fast interrupt 8
  constant trap_firq9_c    : std_ulogic_vector(6 downto 0) := "1" & "0" & "11001"; -- 25: fast interrupt 9
  constant trap_firq10_c   : std_ulogic_vector(6 downto 0) := "1" & "0" & "11010"; -- 26: fast interrupt 10
  constant trap_firq11_c   : std_ulogic_vector(6 downto 0) := "1" & "0" & "11011"; -- 27: fast interrupt 11
  constant trap_firq12_c   : std_ulogic_vector(6 downto 0) := "1" & "0" & "11100"; -- 28: fast interrupt 12
  constant trap_firq13_c   : std_ulogic_vector(6 downto 0) := "1" & "0" & "11101"; -- 29: fast interrupt 13
  constant trap_firq14_c   : std_ulogic_vector(6 downto 0) := "1" & "0" & "11110"; -- 30: fast interrupt 14
  constant trap_firq15_c   : std_ulogic_vector(6 downto 0) := "1" & "0" & "11111"; -- 31: fast interrupt 15
  -- entering debug mode (sync./async. exceptions) --
  constant trap_db_break_c : std_ulogic_vector(6 downto 0) := "0" & "1" & "00001"; -- 1: break instruction (sync)
  constant trap_db_trig_c  : std_ulogic_vector(6 downto 0) := "0" & "1" & "00010"; -- 2: hardware trigger (sync)
  constant trap_db_halt_c  : std_ulogic_vector(6 downto 0) := "1" & "1" & "00011"; -- 3: external halt request (async)
  constant trap_db_step_c  : std_ulogic_vector(6 downto 0) := "1" & "1" & "00100"; -- 4: single-stepping (async)

  -- Trap System ----------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- exception source bits --
  constant exc_iaccess_c  : natural :=  0; -- instruction access fault
  constant exc_illegal_c  : natural :=  1; -- illegal instruction
  constant exc_ialign_c   : natural :=  2; -- instruction address misaligned
  constant exc_ecall_c    : natural :=  3; -- environment call
  constant exc_ebreak_c   : natural :=  4; -- breakpoint
  constant exc_salign_c   : natural :=  5; -- store address misaligned
  constant exc_lalign_c   : natural :=  6; -- load address misaligned
  constant exc_saccess_c  : natural :=  7; -- store access fault
  constant exc_laccess_c  : natural :=  8; -- load access fault
  -- for debug mode only --
  constant exc_db_break_c : natural :=  9; -- enter debug mode via ebreak instruction
  constant exc_db_hw_c    : natural := 10; -- enter debug mode via hw trigger
  --
  constant exc_width_c    : natural := 11; -- length of this list in bits
  -- interrupt source bits --
  constant irq_msi_irq_c  : natural :=  0; -- machine software interrupt
  constant irq_mti_irq_c  : natural :=  1; -- machine timer interrupt
  constant irq_mei_irq_c  : natural :=  2; -- machine external interrupt
  constant irq_firq_0_c   : natural :=  3; -- fast interrupt channel 0
  constant irq_firq_1_c   : natural :=  4; -- fast interrupt channel 1
  constant irq_firq_2_c   : natural :=  5; -- fast interrupt channel 2
  constant irq_firq_3_c   : natural :=  6; -- fast interrupt channel 3
  constant irq_firq_4_c   : natural :=  7; -- fast interrupt channel 4
  constant irq_firq_5_c   : natural :=  8; -- fast interrupt channel 5
  constant irq_firq_6_c   : natural :=  9; -- fast interrupt channel 6
  constant irq_firq_7_c   : natural := 10; -- fast interrupt channel 7
  constant irq_firq_8_c   : natural := 11; -- fast interrupt channel 8
  constant irq_firq_9_c   : natural := 12; -- fast interrupt channel 9
  constant irq_firq_10_c  : natural := 13; -- fast interrupt channel 10
  constant irq_firq_11_c  : natural := 14; -- fast interrupt channel 11
  constant irq_firq_12_c  : natural := 15; -- fast interrupt channel 12
  constant irq_firq_13_c  : natural := 16; -- fast interrupt channel 13
  constant irq_firq_14_c  : natural := 17; -- fast interrupt channel 14
  constant irq_firq_15_c  : natural := 18; -- fast interrupt channel 15
  -- for debug mode only --
  constant irq_db_halt_c  : natural := 19; -- enter debug mode via external halt request
  constant irq_db_step_c  : natural := 20; -- enter debug mode via single-stepping
  --
  constant irq_width_c    : natural := 21; -- length of this list in bits

  -- Privilege Modes ------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant priv_mode_m_c : std_ulogic := '1'; -- machine mode
  constant priv_mode_u_c : std_ulogic := '0'; -- user mode

  -- HPM Event System -----------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  constant hpmcnt_event_cy_c          : natural := 0;  -- Active cycle
  constant hpmcnt_event_tm_c          : natural := 1;  -- Time (unused/reserved)
  constant hpmcnt_event_ir_c          : natural := 2;  -- Retired instruction
  --constant hpmcnt_event_cir_c       : natural := 3;  -- Retired compressed instruction
  --constant hpmcnt_event_wait_if_c   : natural := 4;  -- Instruction fetch memory wait cycle
  --constant hpmcnt_event_wait_ii_c   : natural := 5;  -- Instruction issue wait cycle
  --constant hpmcnt_event_wait_mc_c   : natural := 6;  -- Multi-cycle ALU-operation wait cycle
  --constant hpmcnt_event_load_c      : natural := 7;  -- Load operation
  --constant hpmcnt_event_store_c       : natural := 8;  -- Store operation
  --constant hpmcnt_event_wait_ls_c     : natural := 9;  -- Load/store memory wait cycle
  --constant hpmcnt_event_tbranch_c     : natural := 12; -- Conditional taken branch
  constant hpmcnt_event_ecc_se_imem   : natural := 3; -- Register file single error
  constant hpmcnt_event_ecc_de_imem   : natural := 4; -- Register file double error
  constant hpmcnt_event_ecc_se_dmem   : natural := 5; -- Data memory single error
  constant hpmcnt_event_ecc_de_dmem   : natural := 6; -- Data memory double error
  constant hpmcnt_event_ecc_se_regfile: natural := 7; -- Register file single error
  constant hpmcnt_event_ecc_de_regfile: natural := 8; -- Register file double error
  constant hpmcnt_event_iv            : natural := 9; -- Instruction validator detecting an error
  constant hpmcnt_event_jump_c        : natural := 10; -- Unconditional jump
  constant hpmcnt_event_branch_c      : natural := 11; -- Conditional branch (taken or not taken)
  constant hpmcnt_event_dsp_timeout   : natural := 12; -- One of the DSPs timed out
  constant hpmcnt_event_trap_c        : natural := 13; -- Entered trap
  constant hpmcnt_event_illegal_c     : natural := 14; -- Illegal instruction exception
  --
  constant hpmcnt_event_size_c    : natural := 15; -- length of this list

-- ****************************************************************************************************************************
-- Helper Functions
-- ****************************************************************************************************************************

  function index_size_f(input : natural) return natural;
  function cond_sel_int_f(cond : boolean; val_t : integer; val_f : integer) return integer;
  function cond_sel_natural_f(cond : boolean; val_t : natural; val_f : natural) return natural;
  function cond_sel_suv_f(cond : boolean; val_t : std_ulogic_vector; val_f : std_ulogic_vector) return std_ulogic_vector;
  function cond_sel_string_f(cond : boolean; val_t : string; val_f : string) return string;
  function bool_to_ulogic_f(cond : boolean) return std_ulogic;
  function bin_to_gray_f(input : std_ulogic_vector) return std_ulogic_vector;
  function gray_to_bin_f(input : std_ulogic_vector) return std_ulogic_vector;
  function or_reduce_f(input : std_ulogic_vector) return std_ulogic;
  function and_reduce_f(input : std_ulogic_vector) return std_ulogic;
  function xor_reduce_f(input : std_ulogic_vector) return std_ulogic;
  function su_undefined_f(input : std_ulogic) return boolean;
  function to_hexchar_f(input : std_ulogic_vector(3 downto 0)) return character;
  function to_hstring32_f(input : std_ulogic_vector(31 downto 0)) return string;
  function bit_rev_f(input : std_ulogic_vector) return std_ulogic_vector;
  function is_power_of_two_f(input : natural) return boolean;
  function bswap32_f(input : std_ulogic_vector) return std_ulogic_vector;
  function popcount_f(input : std_ulogic_vector) return natural;
  function leading_zeros_f(input : std_ulogic_vector) return natural;
  impure function mem32_init_f(init : mem32_t; depth : natural) return mem32_t;

-- ****************************************************************************************************************************
-- NEORV32 Processor Top Entity (component prototype)
-- ****************************************************************************************************************************

  component neorv32_top
    generic (
      -- General --
      CLOCK_FREQUENCY            : natural;
      HART_ID                    : std_ulogic_vector(31 downto 0) := x"00000000";
      VENDOR_ID                  : std_ulogic_vector(31 downto 0) := x"00000000";
      INT_BOOTLOADER_EN          : boolean := false;
      -- On-Chip Debugger (OCD) --
      ON_CHIP_DEBUGGER_EN        : boolean := false;
      DM_LEGACY_MODE             : boolean := false;
      -- RISC-V CPU Extensions --
      CPU_EXTENSION_RISCV_A      : boolean := false;
      CPU_EXTENSION_RISCV_B      : boolean := false;
      CPU_EXTENSION_RISCV_C      : boolean := false;
      CPU_EXTENSION_RISCV_E      : boolean := false;
      CPU_EXTENSION_RISCV_M      : boolean := false;
      CPU_EXTENSION_RISCV_U      : boolean := false;
      CPU_EXTENSION_RISCV_Zfinx  : boolean := false;
      CPU_EXTENSION_RISCV_Zicntr : boolean := true;
      CPU_EXTENSION_RISCV_Zihpm  : boolean := false;
      CPU_EXTENSION_RISCV_Zmmul  : boolean := false;
      CPU_EXTENSION_RISCV_Zxcfu  : boolean := false;
      -- Tuning Options --
      FAST_MUL_EN                : boolean := false;
      FAST_SHIFT_EN              : boolean := false;
      REGFILE_HW_RST             : boolean := false;
      -- Physical Memory Protection (PMP) --
      PMP_NUM_REGIONS            : natural range 0 to 16 := 0;
      PMP_MIN_GRANULARITY        : natural := 4;
      -- Hardware Performance Monitors (HPM) --
      HPM_NUM_CNTS               : natural range 0 to 13 := 0;
      HPM_CNT_WIDTH              : natural range 0 to 64 := 40;
      -- Atomic Memory Access - Reservation Set Granularity --
      AMO_RVS_GRANULARITY        : natural := 4;
      -- Internal Instruction memory (IMEM) --
      MEM_INT_IMEM_EN            : boolean := false;
      MEM_INT_IMEM_SIZE          : natural := 16*1024;
      MEM_INT_IMEM_PREFETCH      : boolean := false;
      MEM_INT_PREFETCH_BASE      : std_logic_vector(31 downto 0) := x"00000000";
      MEM_INT_IMEM_SEC           : integer := 1;
      MEM_INT_IV_EN              : boolean := false;
      -- Internal Data memory (DMEM) --
      MEM_INT_DMEM_EN            : boolean := false;
      MEM_INT_DMEM_SIZE          : natural := 8*1024;
      -- Internal Instruction Cache (iCACHE) --
      ICACHE_EN                  : boolean                  := false;
      ICACHE_NUM_BLOCKS          : natural range 1 to 256   := 4;
      ICACHE_BLOCK_SIZE          : natural range 4 to 2**16 := 64;
      ICACHE_ASSOCIATIVITY       : natural range 1 to 2     := 1;
      -- Internal Data Cache (dCACHE) --
      DCACHE_EN                  : boolean                  := false;
      DCACHE_NUM_BLOCKS          : natural range 1 to 256   := 4;
      DCACHE_BLOCK_SIZE          : natural range 4 to 2**16 := 64;
      -- External memory interface (WISHBONE) --
      MEM_EXT_EN                 : boolean := false;
      MEM_EXT_TIMEOUT            : natural := 255;
      MEM_EXT_PIPE_MODE          : boolean := false;
      MEM_EXT_BIG_ENDIAN         : boolean := false;
      MEM_EXT_ASYNC_RX           : boolean := false;
      MEM_EXT_ASYNC_TX           : boolean := false;
      -- External Interrupts Controller (XIRQ) --
      XIRQ_NUM_CH                : natural range 0 to 32          := 0;
      XIRQ_TRIGGER_TYPE          : std_ulogic_vector(31 downto 0) := x"ffffffff";
      XIRQ_TRIGGER_POLARITY      : std_ulogic_vector(31 downto 0) := x"ffffffff";
      -- Processor peripherals --
      IO_GPIO_NUM                : natural range 0 to 64          := 0;
      IO_MTIME_EN                : boolean                        := false;
      IO_UART0_EN                : boolean                        := false;
      IO_UART0_RX_FIFO           : natural range 1 to 2**15       := 1;
      IO_UART0_TX_FIFO           : natural range 1 to 2**15       := 1;
      IO_UART1_EN                : boolean                        := false;
      IO_UART1_RX_FIFO           : natural range 1 to 2**15       := 1;
      IO_UART1_TX_FIFO           : natural range 1 to 2**15       := 1;
      IO_SPI_EN                  : boolean                        := false;
      IO_SPI_FIFO                : natural range 1 to 2**15       := 1;
      IO_SDI_EN                  : boolean                        := false;
      IO_SDI_FIFO                : natural range 1 to 2**15       := 1;
      IO_TWI_EN                  : boolean                        := false;
      IO_PWM_NUM_CH              : natural range 0 to 12          := 0;
      IO_WDT_EN                  : boolean                        := false;
      IO_TRNG_EN                 : boolean                        := false;
      IO_TRNG_FIFO               : natural range 1 to 2**15       := 1;
      IO_CFS_EN                  : boolean                        := false;
      IO_CFS_CONFIG              : std_ulogic_vector(31 downto 0) := x"00000000";
      IO_CFS_IN_SIZE             : natural                        := 32;
      IO_CFS_OUT_SIZE            : natural                        := 32;
      IO_NEOLED_EN               : boolean                        := false;
      IO_NEOLED_TX_FIFO          : natural range 1 to 2**15       := 1;
      IO_GPTMR_EN                : boolean                        := false;
      IO_XIP_EN                  : boolean                        := false;
      IO_ONEWIRE_EN              : boolean                        := false;
      IO_DMA_EN                  : boolean                        := false;
      IO_SLINK_EN                : boolean                        := false;
      IO_SLINK_RX_FIFO           : natural range 1 to 2**15       := 1;
      IO_SLINK_TX_FIFO           : natural range 1 to 2**15       := 1;
      IO_CRC_EN                  : boolean                        := false
    );
    port (
      -- Global control --
      clk_i          : in  std_ulogic;
      rstn_i         : in  std_ulogic;
      -- JTAG on-chip debugger interface --
      jtag_trst_i    : in  std_ulogic := 'U';
      jtag_tck_i     : in  std_ulogic := 'U';
      jtag_tdi_i     : in  std_ulogic := 'U';
      jtag_tdo_o     : out std_ulogic;
      jtag_tms_i     : in  std_ulogic := 'U';
      -- Wishbone bus interface (available if MEM_EXT_EN = true) --
      wb_tag_o       : out std_ulogic_vector(02 downto 0);
      wb_adr_o       : out std_ulogic_vector(31 downto 0);
      wb_dat_i       : in  std_ulogic_vector(31 downto 0) := (others => 'U');
      wb_dat_o       : out std_ulogic_vector(31 downto 0);
      wb_we_o        : out std_ulogic;
      wb_sel_o       : out std_ulogic_vector(03 downto 0);
      wb_stb_o       : out std_ulogic;
      wb_cyc_o       : out std_ulogic;
      wb_ack_i       : in  std_ulogic := 'L';
      wb_err_i       : in  std_ulogic := 'L';
      -- Stream Link Interface (available if IO_SLINK_EN = true) --
      slink_rx_dat_i : in  std_ulogic_vector(31 downto 0) := (others => 'U');
      slink_rx_val_i : in  std_ulogic := 'L';
      slink_rx_rdy_o : out std_ulogic;
      slink_tx_dat_o : out std_ulogic_vector(31 downto 0);
      slink_tx_val_o : out std_ulogic;
      slink_tx_rdy_i : in  std_ulogic := 'L';
      -- Advanced memory control signals --
      fence_o        : out std_ulogic;
      fencei_o       : out std_ulogic;
      -- XIP (execute in place via SPI) signals (available if IO_XIP_EN = true) --
      xip_csn_o      : out std_ulogic;
      xip_clk_o      : out std_ulogic;
      xip_dat_i      : in  std_ulogic := 'L';
      xip_dat_o      : out std_ulogic;
      -- GPIO (available if IO_GPIO_NUM > 0) --
      gpio_o         : out std_ulogic_vector(63 downto 0);
      gpio_i         : in  std_ulogic_vector(63 downto 0) := (others => 'U');
      -- primary UART0 (available if IO_UART0_EN = true) --
      uart0_txd_o    : out std_ulogic;
      uart0_rxd_i    : in  std_ulogic := 'U';
      uart0_rts_o    : out std_ulogic;
      uart0_cts_i    : in  std_ulogic := 'L';
      -- secondary UART1 (available if IO_UART1_EN = true) --
      uart1_txd_o    : out std_ulogic;
      uart1_rxd_i    : in  std_ulogic := 'U'; -- UART1 receive data
      uart1_rts_o    : out std_ulogic;
      uart1_cts_i    : in  std_ulogic := 'L';
      -- SPI (available if IO_SPI_EN = true) --
      spi_clk_o      : out std_ulogic;
      spi_dat_o      : out std_ulogic;
      spi_dat_i      : in  std_ulogic := 'U';
      spi_csn_o      : out std_ulogic_vector(07 downto 0); -- SPI CS
      -- SDI (available if IO_SDI_EN = true) --
      sdi_clk_i      : in  std_ulogic := 'U';
      sdi_dat_o      : out std_ulogic;
      sdi_dat_i      : in  std_ulogic := 'U';
      sdi_csn_i      : in  std_ulogic := 'H';
      -- TWI (available if IO_TWI_EN = true) --
      twi_sda_i      : in  std_ulogic := 'H';
      twi_sda_o      : out std_ulogic;
      twi_scl_i      : in  std_ulogic := 'H';
      twi_scl_o      : out std_ulogic;
      -- 1-Wire Interface (available if IO_ONEWIRE_EN = true) --
      onewire_i      : in  std_ulogic := 'H';
      onewire_o      : out std_ulogic;
      -- PWM (available if IO_PWM_NUM_CH > 0) --
      pwm_o          : out std_ulogic_vector(11 downto 0); -- pwm channels
      -- Custom Functions Subsystem IO --
      cfs_in_i       : in  std_ulogic_vector(IO_CFS_IN_SIZE-1 downto 0) := (others => 'U');
      cfs_out_o      : out std_ulogic_vector(IO_CFS_OUT_SIZE-1 downto 0);
      -- NeoPixel-compatible smart LED interface (available if IO_NEOLED_EN = true) --
      neoled_o       : out std_ulogic;
      -- External platform interrupts (available if XIRQ_NUM_CH > 0) --
      xirq_i         : in  std_ulogic_vector(31 downto 0) := (others => 'L');
      -- CPU Interrupts --
      mtime_irq_i    : in  std_ulogic := 'L';
      msw_irq_i      : in  std_ulogic := 'L';
      mext_irq_i     : in  std_ulogic := 'L'
    );
  end component;

end neorv32_package;

package body neorv32_package is

-- ****************************************************************************************************************************
-- Functions
-- ****************************************************************************************************************************

  -- Minimal required number of bits to represent <input> numbers ---------------------------
  -- -------------------------------------------------------------------------------------------
  function index_size_f(input : natural) return natural is
  begin
    for i in 0 to natural'high loop
      if (2**i >= input) then
        return i;
      end if;
    end loop;
    return 0;
  end function index_size_f;

  -- Conditional select integer -------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function cond_sel_int_f(cond : boolean; val_t : integer; val_f : integer) return integer is
  begin
    if (cond = true) then
      return val_t;
    else
      return val_f;
    end if;
  end function cond_sel_int_f;

  -- Conditional select natural -------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function cond_sel_natural_f(cond : boolean; val_t : natural; val_f : natural) return natural is
  begin
    if (cond = true) then
      return val_t;
    else
      return val_f;
    end if;
  end function cond_sel_natural_f;

  -- Conditional select std_ulogic_vector ---------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function cond_sel_suv_f(cond : boolean; val_t : std_ulogic_vector; val_f : std_ulogic_vector) return std_ulogic_vector is
  begin
    if (cond = true) then
      return val_t;
    else
      return val_f;
    end if;
  end function cond_sel_suv_f;

  -- Conditional select string --------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function cond_sel_string_f(cond : boolean; val_t : string; val_f : string) return string is
  begin
    if (cond = true) then
      return val_t;
    else
      return val_f;
    end if;
  end function cond_sel_string_f;

  -- Convert boolean to std_ulogic ----------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function bool_to_ulogic_f(cond : boolean) return std_ulogic is
  begin
    if (cond = true) then
      return '1';
    else
      return '0';
    end if;
  end function bool_to_ulogic_f;

  -- Convert binary to gray -----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function bin_to_gray_f(input : std_ulogic_vector) return std_ulogic_vector is
    variable tmp_v : std_ulogic_vector(input'range);
  begin
    tmp_v(input'length-1) := input(input'length-1); -- keep MSB
    for i in input'length-2 downto 0 loop
      tmp_v(i) := input(i) xor input(i+1);
    end loop;
    return tmp_v;
  end function bin_to_gray_f;

  -- Convert gray to binary -----------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function gray_to_bin_f(input : std_ulogic_vector) return std_ulogic_vector is
    variable tmp_v : std_ulogic_vector(input'range);
  begin
    tmp_v(input'length-1) := input(input'length-1); -- keep MSB
    for i in input'length-2 downto 0 loop
      tmp_v(i) := tmp_v(i+1) xor input(i);
    end loop;
    return tmp_v;
  end function gray_to_bin_f;

  -- OR all bits ----------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function or_reduce_f(input : std_ulogic_vector) return std_ulogic is
    variable tmp_v : std_ulogic;
  begin
    tmp_v := '0';
    for i in input'range loop
      tmp_v := tmp_v or input(i);
    end loop;
    return tmp_v;
  end function or_reduce_f;

  -- AND all bits ---------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function and_reduce_f(input : std_ulogic_vector) return std_ulogic is
    variable tmp_v : std_ulogic;
  begin
    tmp_v := '1';
    for i in input'range loop
      tmp_v := tmp_v and input(i);
    end loop;
    return tmp_v;
  end function and_reduce_f;

  -- XOR all bits ---------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function xor_reduce_f(input : std_ulogic_vector) return std_ulogic is
    variable tmp_v : std_ulogic;
  begin
    tmp_v := '0';
    for i in input'range loop
      tmp_v := tmp_v xor input(i);
    end loop;
    return tmp_v;
  end function xor_reduce_f;

  -- Check if std_ulogic is not '1' or '0' --------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function su_undefined_f(input : std_ulogic) return boolean is
  begin
    case input is
      when '1' | '0' => return false;
      when others    => return true;
    end case;
  end function su_undefined_f;

  -- Convert std_ulogic_vector to lowercase HEX char ----------------------------------------
  -- -------------------------------------------------------------------------------------------
  function to_hexchar_f(input : std_ulogic_vector(3 downto 0)) return character is
    variable hex_v : string(1 to 16);
  begin
    hex_v := "0123456789abcdef";
    if (su_undefined_f(input(3)) = true) or (su_undefined_f(input(2)) = true) or
       (su_undefined_f(input(1)) = true) or (su_undefined_f(input(0)) = true) then
      return '?';
    else
      return hex_v(to_integer(unsigned(input)) + 1);
    end if;
  end function to_hexchar_f;

  -- Convert 32-bit std_ulogic_vector to hex string -----------------------------------------
  -- -------------------------------------------------------------------------------------------
  function to_hstring32_f(input : std_ulogic_vector(31 downto 0)) return string is
    variable res_v : string(1 to 8);
  begin
    for i in 7 downto 0 loop
      res_v(8-i) := to_hexchar_f(input(i*4+3 downto i*4+0));
    end loop;
    return res_v;
  end function to_hstring32_f;

  -- Bit reversal ---------------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function bit_rev_f(input : std_ulogic_vector) return std_ulogic_vector is
    variable output_v : std_ulogic_vector(input'range);
  begin
    for i in 0 to input'length-1 loop
      output_v(input'length-i-1) := input(i);
    end loop;
    return output_v;
  end function bit_rev_f;

  -- Test if input number is a power of two -------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function is_power_of_two_f(input : natural) return boolean is
    variable tmp : unsigned(31 downto 0);
  begin
    if (input = 0) then
      return false;
    elsif (input = 1) then
      return true;
    else
      tmp := to_unsigned(input, 32);
      if ((tmp and (tmp - 1)) = 0) then
        return true;
      else
        return false;
      end if;
    end if;
  end function is_power_of_two_f;

  -- Swap all bytes of a 32-bit word (endianness conversion) --------------------------------
  -- -------------------------------------------------------------------------------------------
  function bswap32_f(input : std_ulogic_vector) return std_ulogic_vector is
    variable output_v : std_ulogic_vector(input'range);
  begin
    output_v(07 downto 00) := input(31 downto 24);
    output_v(15 downto 08) := input(23 downto 16);
    output_v(23 downto 16) := input(15 downto 08);
    output_v(31 downto 24) := input(07 downto 00);
    return output_v;
  end function bswap32_f;

  -- Population count (number of set bits) --------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function popcount_f(input : std_ulogic_vector) return natural is
    variable cnt_v : natural range 0 to input'length;
  begin
    cnt_v := 0;
    for i in input'length-1 downto 0 loop
      if (input(i) = '1') then
        cnt_v := cnt_v + 1;
      end if;
    end loop;
    return cnt_v;
  end function popcount_f;

  -- Count leading zeros --------------------------------------------------------------------
  -- -------------------------------------------------------------------------------------------
  function leading_zeros_f(input : std_ulogic_vector) return natural is
    variable cnt_v : natural range 0 to input'length;
  begin
    cnt_v := 0;
    for i in input'length-1 downto 0 loop
      if (input(i) = '0') then
        cnt_v := cnt_v + 1;
      else
        exit;
      end if;
    end loop;
    return cnt_v;
  end function leading_zeros_f;

  -- Initialize mem32_t array from another mem32_t array ------------------------------------
  -- -------------------------------------------------------------------------------------------
  impure function mem32_init_f(init : mem32_t; depth : natural) return mem32_t is
    variable mem_v : mem32_t(0 to depth-1);
  begin
    mem_v := (others => (others => '0')); -- [IMPORTANT] make sure remaining memory entries are set to zero
    if (init'length > depth) then
      return mem_v;
    end if;
    for i in 0 to init'length-1 loop -- initialize only in range of source data array
      mem_v(i) := init(i);
    end loop;
    return mem_v;
  end function mem32_init_f;


end neorv32_package;

-- ****************************************************************************************************************************
-- Additional Packages
-- ****************************************************************************************************************************

  -- Prototype Definition: bootloader_init_image --------------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- > memory content in 'neorv32_bootloader_image.vhd', auto-generated by 'image_gen'
  -- > used by 'neorv32_boot_rom.vhd'
  -- > enables body-only recompile in case of firmware change (NEORV32 PR #338)

library ieee;
use ieee.std_logic_1164.all;

library neorv32;
use neorv32.neorv32_package.all;

package neorv32_bootloader_image is
  constant bootloader_init_image : mem32_t;
end neorv32_bootloader_image;


  -- Prototype Definition: neorv32_application_image ----------------------------------------
  -- -------------------------------------------------------------------------------------------
  -- > memory content in 'neorv32_application_image.vhd', auto-generated by 'image_gen'
  -- > used by 'mem/neorv32_imem.*.vhd'
  -- > enables body-only recompile in case of firmware change (NEORV32 PR #338)

library ieee;
use ieee.std_logic_1164.all;

library neorv32;
use neorv32.neorv32_package.all;

package neorv32_application_image is
  constant application_init_image : mem32_t := (
x"de067139",
x"0080dc22",
x"fca42623",
x"152387ae",
x"1723fcf4",
x"1623fe04",
x"1523fe04",
x"2783fe04",
x"53dcfcc4",
x"fef42223",
x"fcc42783",
x"0047d783",
x"fcf41e23",
x"fca45783",
x"fcf41923",
x"fc041f23",
x"5783a221",
x"f793fde4",
x"07c20ff7",
x"182387c1",
x"0793fcf4",
x"85befd04",
x"fe442503",
x"2a232ad5",
x"2503fca4",
x"24b5fe44",
x"fea42223",
x"fd442783",
x"5783eb95",
x"0785fea4",
x"fef41523",
x"fe442783",
x"43dc439c",
x"00079783",
x"07c287a1",
x"07c287c1",
x"8b8583c1",
x"83c107c2",
x"fee45703",
x"172397ba",
x"a89dfef4",
x"fec45783",
x"16230785",
x"2783fef4",
x"43dcfd44",
x"00079783",
x"83c107c2",
x"c39d8b85",
x"fd442783",
x"978343dc",
x"87a50007",
x"87c107c2",
x"83c107c2",
x"07c28b85",
x"570383c1",
x"97bafee4",
x"fef41723",
x"fd442783",
x"c79d439c",
x"fd442783",
x"2023439c",
x"2783fef4",
x"4398fe04",
x"fd442783",
x"2783c398",
x"4398fe44",
x"fe042783",
x"2783c398",
x"2703fe44",
x"c398fe04",
x"fd241783",
x"0007cd63",
x"fd241783",
x"83c107c2",
x"07c20785",
x"07c283c1",
x"192387c1",
x"1783fcf4",
x"07c2fde4",
x"078583c1",
x"83c107c2",
x"fcf41f23",
x"fde41703",
x"fdc41783",
x"eef749e3",
x"fec45783",
x"07c2078a",
x"570383c1",
x"8f99fea4",
x"83c107c2",
x"fee45703",
x"172397ba",
x"1783fef4",
x"5b63fca4",
x"260300f0",
x"0593fcc4",
x"25035660",
x"2c25fe44",
x"fea42223",
x"fe442783",
x"853e439c",
x"2c232251",
x"0793fca4",
x"85befd04",
x"fe442503",
x"20232075",
x"2783fea4",
x"eb95fe04",
x"fe442783",
x"2023439c",
x"a025fef4",
x"fe442783",
x"978343dc",
x"57030007",
x"85bafee4",
x"00ef853e",
x"87aa4050",
x"fef41723",
x"fe042783",
x"2023439c",
x"2783fef4",
x"fbf9fe04",
x"fe442783",
x"85be439c",
x"fd842503",
x"2c232aad",
x"4601fca4",
x"5b400593",
x"fe442503",
x"22232a6d",
x"2783fea4",
x"439cfe44",
x"fef42023",
x"2783a025",
x"43dcfe44",
x"00079783",
x"fee45703",
x"853e85ba",
x"3ab000ef",
x"172387aa",
x"2783fef4",
x"439cfe04",
x"fef42023",
x"fe042783",
x"5783fbf9",
x"853efee4",
x"546250f2",
x"80826121",
x"ce221101",
x"26231000",
x"2423fea4",
x"2783feb4",
x"9783fe84",
x"ce630027",
x"a0310207",
x"fec42783",
x"2623439c",
x"2783fef4",
x"cf81fec4",
x"fec42783",
x"970343dc",
x"27830027",
x"9783fe84",
x"1fe30027",
x"2783fcf7",
x"a815fec4",
x"fec42783",
x"2623439c",
x"2783fef4",
x"c385fec4",
x"fec42783",
x"978343dc",
x"07c20007",
x"f79383c1",
x"27030ff7",
x"1703fe84",
x"9be30007",
x"2783fce7",
x"853efec4",
x"61054472",
x"71798082",
x"1800d622",
x"fca42e23",
x"fe042623",
x"2783a01d",
x"439cfdc4",
x"fef42423",
x"fdc42783",
x"fec42703",
x"2783c398",
x"2623fdc4",
x"2783fef4",
x"2e23fe84",
x"2783fcf4",
x"ffe1fdc4",
x"fec42783",
x"5432853e",
x"80826145",
x"d6227179",
x"2e231800",
x"2783fca4",
x"439cfdc4",
x"fef42623",
x"fdc42783",
x"242343dc",
x"2783fef4",
x"43d8fec4",
x"fdc42783",
x"2783c3d8",
x"2703fec4",
x"c3d8fe84",
x"fdc42783",
x"4398439c",
x"fdc42783",
x"2783c398",
x"a023fec4",
x"27830007",
x"853efec4",
x"61455432",
x"71798082",
x"1800d622",
x"fca42e23",
x"fcb42c23",
x"fdc42783",
x"262343dc",
x"2783fef4",
x"43d8fd84",
x"fdc42783",
x"2783c3d8",
x"2703fd84",
x"c3d8fec4",
x"fd842783",
x"27834398",
x"c398fdc4",
x"fd842783",
x"fdc42703",
x"2783c398",
x"853efdc4",
x"61455432",
x"715d8082",
x"c4a2c686",
x"2e230880",
x"2c23faa4",
x"2a23fab4",
x"4785fac4",
x"fcf42e23",
x"fbc42783",
x"fef42623",
x"fa042e23",
x"fe042023",
x"fc042c23",
x"2783a291",
x"0785fd84",
x"fcf42c23",
x"fec42783",
x"fef42423",
x"fc042a23",
x"fc042623",
x"2783a01d",
x"0785fd44",
x"fcf42a23",
x"fe842783",
x"2423439c",
x"2783fef4",
x"cf89fe84",
x"fcc42783",
x"26230785",
x"2703fcf4",
x"2783fcc4",
x"4ae3fdc4",
x"a011fcf7",
x"27830001",
x"2823fdc4",
x"a0f1fcf4",
x"fd442783",
x"2783e385",
x"2223fe84",
x"2783fef4",
x"439cfe84",
x"fef42423",
x"fd042783",
x"282317fd",
x"a059fcf4",
x"fd042783",
x"2783c781",
x"e385fe84",
x"fec42783",
x"fef42223",
x"fec42783",
x"2623439c",
x"2783fef4",
x"17fdfd44",
x"fcf42a23",
x"2783a8b1",
x"43d8fec4",
x"fe842783",
x"278343d4",
x"2603fb84",
x"85b6fb44",
x"9782853a",
x"416387aa",
x"278302f0",
x"2223fec4",
x"2783fef4",
x"439cfec4",
x"fef42623",
x"fd442783",
x"2a2317fd",
x"a839fcf4",
x"fe842783",
x"fef42223",
x"fe842783",
x"2423439c",
x"2783fef4",
x"17fdfd04",
x"fcf42823",
x"fe042783",
x"2783c799",
x"2703fe04",
x"c398fe44",
x"2783a029",
x"2e23fe44",
x"2783faf4",
x"2023fe44",
x"2783fef4",
x"49e3fd44",
x"2783f2f0",
x"5563fd04",
x"278300f0",
x"f38dfe84",
x"fe842783",
x"fef42623",
x"fec42783",
x"ea079de3",
x"fe042783",
x"0007a023",
x"fd842703",
x"c5634785",
x"278300e7",
x"a039fbc4",
x"fdc42783",
x"2e230786",
x"bdbdfcf4",
x"40b6853e",
x"61614426",
x"71798082",
x"d422d606",
x"2e231800",
x"2c23fca4",
x"2a23fcb4",
x"2783fcc4",
x"2583fdc4",
x"853efd44",
x"87aa28d9",
x"fef41723",
x"fd842783",
x"fd442583",
x"20d1853e",
x"162387aa",
x"1703fef4",
x"1783fee4",
x"07b3fec4",
x"853e40f7",
x"542250b2",
x"80826145",
x"ce221101",
x"26231000",
x"2423fea4",
x"2223feb4",
x"2783fec4",
x"ebadfe44",
x"fec42783",
x"00079783",
x"f007f793",
x"01079713",
x"27838741",
x"9783fec4",
x"07c20007",
x"83a183c1",
x"83c107c2",
x"87c107c2",
x"97138fd9",
x"87410107",
x"fec42783",
x"00e79023",
x"fe842783",
x"00079783",
x"f007f793",
x"01079713",
x"27838741",
x"9783fe84",
x"07c20007",
x"83a183c1",
x"83c107c2",
x"87c107c2",
x"97138fd9",
x"87410107",
x"fe842783",
x"00e79023",
x"fec42783",
x"00279783",
x"2783873e",
x"9783fe84",
x"07b30027",
x"853e40f7",
x"61054472",
x"71798082",
x"d422d606",
x"2e231800",
x"2c23fca4",
x"2783fcb4",
x"d783fdc4",
x"15230007",
x"1783fef4",
x"879dfea4",
x"87c107c2",
x"0ff7f793",
x"04a38b85",
x"4783fef4",
x"cb81fe94",
x"fea45783",
x"07f7f793",
x"87c107c2",
x"5783aa2d",
x"8b9dfea4",
x"fef41323",
x"fea41783",
x"07c2878d",
x"8bbd87c1",
x"fef41623",
x"fec45783",
x"07c20792",
x"570387c1",
x"8fd9fec4",
x"fef41623",
x"fe641783",
x"4705c789",
x"06e78163",
x"1703a861",
x"0793fec4",
x"c6630210",
x"079300e7",
x"16230220",
x"2783fef4",
x"4f88fd84",
x"fd842783",
x"27834bcc",
x"9603fd84",
x"27830007",
x"9683fd84",
x"27830027",
x"d783fd84",
x"17030387",
x"26c5fec4",
x"172387aa",
x"2783fef4",
x"d783fd84",
x"ebb103e7",
x"fee45703",
x"fd842783",
x"02e79f23",
x"2783a099",
x"8713fd84",
x"27830287",
x"d683fd84",
x"17830387",
x"8636fec4",
x"853a85be",
x"87aa2605",
x"fef41723",
x"fd842783",
x"03c7d783",
x"5703ef99",
x"2783fee4",
x"9e23fd84",
x"a80102e7",
x"fea45783",
x"fef41723",
x"0001a021",
x"0001a011",
x"fee45703",
x"fd842783",
x"0387d783",
x"853a85be",
x"87aa2d8d",
x"2783873e",
x"9c23fd84",
x"578302e7",
x"f793fee4",
x"172307f7",
x"5783fef4",
x"f793fea4",
x"07c2f007",
x"e79387c1",
x"07c20807",
x"570387c1",
x"8fd9fee4",
x"01079713",
x"27838741",
x"9023fdc4",
x"178300e7",
x"853efee4",
x"542250b2",
x"80826145",
x"d6067179",
x"1800d422",
x"fca42e23",
x"fdc42783",
x"fef42423",
x"fe842783",
x"22234fdc",
x"2783fef4",
x"9c23fe84",
x"27830207",
x"9d23fe84",
x"27830207",
x"9e23fe84",
x"27830207",
x"9f23fe84",
x"26230207",
x"a8bdfe04",
x"25034585",
x"f0effe84",
x"87aafd6f",
x"fef41123",
x"fe842783",
x"0387d703",
x"fe245783",
x"853e85ba",
x"87aa2b7d",
x"2783873e",
x"9c23fe84",
x"55fd02e7",
x"fe842503",
x"fa8ff0ef",
x"112387aa",
x"2783fef4",
x"d703fe84",
x"57830387",
x"85bafe24",
x"2b41853e",
x"873e87aa",
x"fe842783",
x"02e79c23",
x"fec42783",
x"2783eb89",
x"d703fe84",
x"27830387",
x"9d23fe84",
x"278302e7",
x"0785fec4",
x"fef42623",
x"fec42703",
x"fe442783",
x"f6f76ee3",
x"853e4781",
x"542250b2",
x"80826145",
x"de227139",
x"26230080",
x"2423fca4",
x"2223fcb4",
x"2023fcc4",
x"2023fcd4",
x"4785fe04",
x"fef42623",
x"fe042423",
x"fe042223",
x"fc442783",
x"4785e38d",
x"fcf42223",
x"2783a829",
x"0785fe84",
x"fef42423",
x"fe842783",
x"02f787b3",
x"2223078e",
x"2703fef4",
x"2783fe44",
x"60e3fcc4",
x"2783fef7",
x"17fdfe84",
x"fef42023",
x"fc842783",
x"9bf117fd",
x"2e230791",
x"2783fcf4",
x"87b3fe04",
x"078602f7",
x"fdc42703",
x"2c2397ba",
x"2423fcf4",
x"a8e9fe04",
x"fe042223",
x"2703a87d",
x"2783fec4",
x"0733fc44",
x"579302f7",
x"83c141f7",
x"00f706b3",
x"177d6741",
x"07b38f75",
x"222340f7",
x"2783fcf4",
x"9713fc44",
x"83410107",
x"fec42783",
x"83c107c2",
x"07c297ba",
x"1b2383c1",
x"2703fcf4",
x"2783fe84",
x"0733fe04",
x"278302f7",
x"97bafe44",
x"27030786",
x"97bafd84",
x"fd645703",
x"00e79023",
x"fec42783",
x"01079713",
x"57838341",
x"97bafd64",
x"83c107c2",
x"fcf41b23",
x"fd645783",
x"0ff7f793",
x"fcf41b23",
x"fe842703",
x"fe042783",
x"02f70733",
x"fe442783",
x"078697ba",
x"fdc42703",
x"570397ba",
x"9023fd64",
x"278300e7",
x"0785fec4",
x"fef42623",
x"fe442783",
x"22230785",
x"2703fef4",
x"2783fe44",
x"6ee3fe04",
x"2783f2f7",
x"0785fe84",
x"fef42423",
x"fe842703",
x"fe042783",
x"f2f760e3",
x"fc042783",
x"fdc42703",
x"2783c3d8",
x"2703fc04",
x"c798fd84",
x"fe042783",
x"02f787b3",
x"27030786",
x"97bafd84",
x"9bf117fd",
x"873e0791",
x"fc042783",
x"2703c7d8",
x"2783fe04",
x"c398fc04",
x"fe042783",
x"5472853e",
x"80826121",
x"de067139",
x"0080dc22",
x"fca42623",
x"873287ae",
x"fcf41523",
x"142387ba",
x"2783fcf4",
x"439cfcc4",
x"fef42623",
x"fcc42783",
x"242347dc",
x"2783fef4",
x"43dcfcc4",
x"fef42223",
x"fcc42783",
x"2023479c",
x"5783fef4",
x"1f23fca4",
x"1783fcf4",
x"873efde4",
x"fe042683",
x"fe442603",
x"fe842583",
x"fec42503",
x"448090ef",
x"873e87aa",
x"fc845783",
x"853a85be",
x"87aa2ccd",
x"fcf41423",
x"fc845783",
x"50f2853e",
x"61215462",
x"71598082",
x"d4a2d686",
x"2e231880",
x"2c23f8a4",
x"85b2f8b4",
x"86ba8636",
x"87ae873e",
x"f8f41b23",
x"1a2387b2",
x"87b6f8f4",
x"f8f41923",
x"182387ba",
x"2783f8f4",
x"2023f984",
x"2623faf4",
x"a81dfe04",
x"fec42783",
x"17c1078a",
x"aa2397a2",
x"2783fa07",
x"078afec4",
x"97a217c1",
x"fb47a703",
x"fec42783",
x"17c1078a",
x"aa2397a2",
x"2783fce7",
x"0785fec4",
x"fef42623",
x"fec42703",
x"f3e3479d",
x"a81dfce7",
x"fa440713",
x"fa040793",
x"853e85ba",
x"3860a0ef",
x"fea42223",
x"fe442783",
x"17c1078a",
x"a78397a2",
x"8713fd47",
x"27830017",
x"078afe44",
x"97a217c1",
x"fce7aa23",
x"fa042783",
x"0007c783",
x"2783f3f1",
x"2023f984",
x"a83dfaf4",
x"fa042783",
x"0007c703",
x"02c00793",
x"02f70163",
x"fa042783",
x"0007c683",
x"f9645783",
x"0ff7f713",
x"fa042783",
x"77138f35",
x"80230ff7",
x"270300e7",
x"1783fa04",
x"97baf924",
x"faf42023",
x"f9842703",
x"f9c42783",
x"2783973e",
x"ebe3fa04",
x"2783fae7",
x"2023f984",
x"a81dfaf4",
x"fa440713",
x"fa040793",
x"853e85ba",
x"2e60a0ef",
x"fea42423",
x"fe842783",
x"17c1078a",
x"a78397a2",
x"8713fd47",
x"27830017",
x"078afe84",
x"97a217c1",
x"fce7aa23",
x"fa042783",
x"0007c783",
x"2783f3f1",
x"2023f984",
x"a83dfaf4",
x"fa042783",
x"0007c703",
x"02c00793",
x"02f70163",
x"fa042783",
x"0007c683",
x"f9445783",
x"0ff7f713",
x"fa042783",
x"77138f35",
x"80230ff7",
x"270300e7",
x"1783fa04",
x"97baf924",
x"faf42023",
x"f9842703",
x"f9c42783",
x"2783973e",
x"ebe3fa04",
x"2623fae7",
x"a0a1fe04",
x"fec42783",
x"17c1078a",
x"a78397a2",
x"5703fd47",
x"85baf904",
x"2a59853e",
x"182387aa",
x"2783f8f4",
x"078afec4",
x"97a217c1",
x"fb47a783",
x"f9045703",
x"853e85ba",
x"87aa2aa5",
x"f8f41823",
x"fec42783",
x"26230785",
x"2703fef4",
x"479dfec4",
x"fae7fae3",
x"f9045783",
x"50b6853e",
x"61655426",
x"71798082",
x"1800d622",
x"872e87aa",
x"fcf40fa3",
x"1e2387ba",
x"07a3fcf4",
x"06a3fe04",
x"0723fe04",
x"07a3fe04",
x"a069fe04",
x"fdc45783",
x"01879713",
x"07838761",
x"8fb9fdf4",
x"87e107e2",
x"0ff7f793",
x"06a38b85",
x"4783fef4",
x"8385fdf4",
x"fcf40fa3",
x"fed44703",
x"1e634785",
x"578300f7",
x"873efdc4",
x"07896791",
x"1e238fb9",
x"4785fcf4",
x"fef40723",
x"0723a019",
x"5783fe04",
x"8385fdc4",
x"fcf41e23",
x"fee44783",
x"5783cb89",
x"873efdc4",
x"8fd977e1",
x"fcf41e23",
x"5783a809",
x"873efdc4",
x"17fd67a1",
x"1e238ff9",
x"4783fcf4",
x"0785fef4",
x"fef407a3",
x"fef44703",
x"f9e3479d",
x"5783f6e7",
x"853efdc4",
x"61455432",
x"11018082",
x"cc22ce06",
x"87aa1000",
x"1723872e",
x"87bafef4",
x"fef41623",
x"fee45783",
x"fec45703",
x"853e85ba",
x"87aa2039",
x"40f2853e",
x"61054462",
x"11018082",
x"cc22ce06",
x"87aa1000",
x"1723872e",
x"87bafef4",
x"fef41623",
x"fee45783",
x"0ff7f793",
x"fec45703",
x"853e85ba",
x"87aa35dd",
x"fef41623",
x"fee45783",
x"07c283a1",
x"f79383c1",
x"57030ff7",
x"85bafec4",
x"35e1853e",
x"162387aa",
x"5783fef4",
x"853efec4",
x"446240f2",
x"80826105",
x"ce061101",
x"1000cc22",
x"fea42623",
x"152387ae",
x"2783fef4",
x"07c2fec4",
x"570387c1",
x"85bafea4",
x"3f91853e",
x"152387aa",
x"2783fef4",
x"83c1fec4",
x"87c107c2",
x"fea45703",
x"853e85ba",
x"87aa3f2d",
x"fef41523",
x"fea45783",
x"40f2853e",
x"61054462",
x"00008082",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"7fff9197",
x"86818193",
x"00000013",
x"00000013",
x"48818113",
x"ff017113",
x"00000297",
x"12028293",
x"30529073",
x"00000097",
x"0a608093",
x"00008563",
x"00ef9082",
x"25730240",
x"4581f140",
x"30ef4601",
x"02977850",
x"82930000",
x"907300c2",
x"23033052",
x"bff50000",
x"42970000",
x"82930000",
x"8317fda2",
x"03137fff",
x"8397fa23",
x"83937fff",
x"8c630163",
x"5a630062",
x"a5030073",
x"02910002",
x"00a32023",
x"4ae30311",
x"8082fe73",
x"b37346a1",
x"42913006",
x"0055c563",
x"00357613",
x"0023ca11",
x"05050005",
x"47e315fd",
x"1073feb0",
x"80823003",
x"00052023",
x"15f10511",
x"fcb04ee3",
x"30031073",
x"20238082",
x"03110003",
x"fe734de3",
x"84068082",
x"ffff8297",
x"f3528293",
x"04028163",
x"ffff8297",
x"f2828293",
x"f14027f3",
x"b07346a1",
x"830a3006",
x"ffff8397",
x"31438393",
x"0363938a",
x"37d10073",
x"00579d63",
x"7fff8317",
x"f0030313",
x"7fff8397",
x"f7438393",
x"00730363",
x"8317376d",
x"03137fff",
x"8397f6a3",
x"83937fff",
x"57637d23",
x"20230073",
x"03110003",
x"fe734de3",
x"808280a2",
x"342022f3",
x"34102373",
x"343023f3",
x"0000bfd5",
x"74617453",
x"00006369",
x"70616548",
x"00000000",
x"63617453",
x"0000006b",
x"65726f43",
x"6b72614d",
x"7a695320",
x"20202065",
x"25203a20",
x"000a756c",
x"61746f54",
x"6974206c",
x"20736b63",
x"20202020",
x"25203a20",
x"6b20756c",
x"0000000a",
x"61746f54",
x"6974206c",
x"2820656d",
x"73636573",
x"25203a29",
x"00000a64",
x"72657449",
x"6f697461",
x"532f736e",
x"20206365",
x"25203a20",
x"00000a64",
x"4f525245",
x"4d202152",
x"20747375",
x"63657865",
x"20657475",
x"20726f66",
x"6c207461",
x"74736165",
x"20303120",
x"73636573",
x"726f6620",
x"76206120",
x"64696c61",
x"73657220",
x"21746c75",
x"0000000a",
x"72657449",
x"6f697461",
x"2020736e",
x"20202020",
x"25203a20",
x"000a756c",
x"31434347",
x"2e322e33",
x"00000030",
x"706d6f43",
x"72656c69",
x"72657620",
x"6e6f6973",
x"25203a20",
x"00000a73",
x"64203e2d",
x"75616665",
x"202c746c",
x"20656573",
x"656b616d",
x"656c6966",
x"00000000",
x"706d6f43",
x"72656c69",
x"616c6620",
x"20207367",
x"25203a20",
x"00000a73",
x"54415453",
x"00004349",
x"6f6d654d",
x"6c207972",
x"7461636f",
x"206e6f69",
x"25203a20",
x"00000a73",
x"64656573",
x"20637263",
x"20202020",
x"20202020",
x"30203a20",
x"34302578",
x"00000a78",
x"5d64255b",
x"6c637263",
x"20747369",
x"20202020",
x"203a2020",
x"30257830",
x"000a7834",
x"5d64255b",
x"6d637263",
x"69727461",
x"20202078",
x"203a2020",
x"30257830",
x"000a7834",
x"5d64255b",
x"73637263",
x"65746174",
x"20202020",
x"203a2020",
x"30257830",
x"000a7834",
x"5d64255b",
x"66637263",
x"6c616e69",
x"20202020",
x"203a2020",
x"30257830",
x"000a7834",
x"72726f43",
x"20746365",
x"7265706f",
x"6f697461",
x"6176206e",
x"6164696c",
x"2e646574",
x"65655320",
x"41455220",
x"2e454d44",
x"6620646d",
x"7220726f",
x"61206e75",
x"7220646e",
x"726f7065",
x"676e6974",
x"6c757220",
x"0a2e7365",
x"00000000",
x"6f727245",
x"64207372",
x"63657465",
x"0a646574",
x"00000000",
x"6e6e6143",
x"7620746f",
x"64696c61",
x"20657461",
x"7265706f",
x"6f697461",
x"6f66206e",
x"68742072",
x"20657365",
x"64656573",
x"6c617620",
x"2c736575",
x"656c7020",
x"20657361",
x"706d6f63",
x"20657261",
x"68746977",
x"73657220",
x"73746c75",
x"206e6f20",
x"6e6b2061",
x"206e776f",
x"74616c70",
x"6d726f66",
x"00000a2e",
x"4f454e0a",
x"32335652",
x"6148203a",
x"61776472",
x"50206572",
x"6f667265",
x"6e616d72",
x"4d206563",
x"74696e6f",
x"2073726f",
x"776f6c28",
x"726f7720",
x"6f207364",
x"29796c6e",
x"0000000a",
x"32313035",
x"00000000",
x"34333231",
x"00000000",
x"3437382d",
x"00000000",
x"3232312b",
x"00000000",
x"352e3533",
x"30303434",
x"00000000",
x"3332312e",
x"30303534",
x"00000000",
x"3031312d",
x"3030372e",
x"00000000",
x"362e302b",
x"30303434",
x"00000000",
x"30352e35",
x"332b6530",
x"00000000",
x"32312e2d",
x"322d6533",
x"00000000",
x"6537382d",
x"3233382b",
x"00000000",
x"362e302b",
x"32312d65",
x"00000000",
x"332e3054",
x"46312d65",
x"00000000",
x"542e542d",
x"71542b2b",
x"00000000",
x"2e335431",
x"7a346534",
x"00000000",
x"302e3433",
x"5e542d65",
x"00000000",
x"0000af68",
x"0000b14a",
x"0000afd4",
x"0000b0b6",
x"0000b028",
x"0000b06a",
x"0000b0f6",
x"0000b12a",
x"0000b1f0",
x"0000b1b6",
x"0000b1c0",
x"0000b1ca",
x"0000b1d8",
x"0000b1e6",
x"4f525245",
x"50203a52",
x"7361656c",
x"6f6d2065",
x"79666964",
x"65687420",
x"74616420",
x"70797461",
x"69207365",
x"6f63206e",
x"705f6572",
x"6d74726f",
x"21682e65",
x"0000000a",
x"33323130",
x"37363534",
x"62613938",
x"66656463",
x"6a696867",
x"6e6d6c6b",
x"7271706f",
x"76757473",
x"7a797877",
x"00000000",
x"33323130",
x"37363534",
x"42413938",
x"46454443",
x"4a494847",
x"4e4d4c4b",
x"5251504f",
x"56555453",
x"5a595857",
x"00000000",
x"4c554e3c",
x"00003e4c",
x"0000b9f6",
x"0000ba20",
x"0000ba20",
x"0000ba04",
x"0000ba20",
x"0000ba20",
x"0000ba20",
x"0000ba20",
x"0000ba20",
x"0000ba20",
x"0000ba20",
x"0000b9e8",
x"0000ba20",
x"0000b9da",
x"0000ba20",
x"0000ba20",
x"0000ba12",
x"0000bd24",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bd96",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bd30",
x"0000bdb8",
x"0000bb90",
x"0000bdaa",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdaa",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bdb8",
x"0000bd8e",
x"0000bcdc",
x"0000bdb8",
x"0000bdb8",
x"0000bc0c",
x"0000bdb8",
x"0000be0c",
x"0000bdb8",
x"0000bdb8",
x"0000bda2",
x"74696e49",
x"6d6f6320",
x"74656c70",
x"000a0d65",
x"ce221101",
x"26231000",
x"0793fea4",
x"439ce000",
x"4472853e",
x"80826105",
x"c6221141",
x"07930800",
x"4798e000",
x"8ff967a1",
x"4785c399",
x"4781a011",
x"4432853e",
x"80820141",
x"c6061141",
x"0800c422",
x"87aa3fe1",
x"40b2853e",
x"01414422",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"30579073",
x"44720001",
x"80826105",
x"ce221101",
x"27f31000",
x"26233420",
x"2783fef4",
x"853efec4",
x"61054472",
x"71798082",
x"d422d606",
x"2e231800",
x"2783fca4",
x"9bf1fdc4",
x"fef42623",
x"fec42503",
x"00013f4d",
x"542250b2",
x"80826145",
x"00000000",
x"00000000",
x"00000000",
x"ce86711d",
x"ca9acc96",
x"c6a2c89e",
x"c2aec4aa",
x"de36c0b2",
x"da3edc3a",
x"d646d842",
x"d276d472",
x"ce7ed07a",
x"37791080",
x"faa42623",
x"fac42783",
x"242383fd",
x"2783faf4",
x"f793fac4",
x"22233ff7",
x"2703faf4",
x"4785fa84",
x"00f71d63",
x"800007b7",
x"0a078713",
x"fa442783",
x"97ba078a",
x"9782439c",
x"8713a819",
x"27838781",
x"078afa44",
x"439c97ba",
x"fa442503",
x"00019782",
x"42e640f6",
x"43c64356",
x"45264436",
x"46064596",
x"576256f2",
x"584257d2",
x"5e2258b2",
x"5f025e92",
x"61254ff2",
x"30200073",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"00000000",
x"ce061101",
x"1000cc22",
x"fe042623",
x"8713a005",
x"27838781",
x"078afec4",
x"672197ba",
x"13870713",
x"2783c398",
x"0785fec4",
x"fef42623",
x"fec42703",
x"fee347bd",
x"67a1fce7",
x"78078513",
x"00013d69",
x"446240f2",
x"80826105",
x"c6061141",
x"0800c422",
x"00013f45",
x"442240b2",
x"80820141",
x"ce221101",
x"87aa1000",
x"fef407a3",
x"77fd0001",
x"50078793",
x"07b74398",
x"8ff90020",
x"77fdfbed",
x"50078793",
x"fef44703",
x"0001c3d8",
x"61054472",
x"71798082",
x"d422d606",
x"2e231800",
x"2c23fca4",
x"20c1fcb4",
x"cbcd87aa",
x"fe042623",
x"fe042423",
x"879377fd",
x"a0235007",
x"27830007",
x"0786fd84",
x"fdc42703",
x"02f757b3",
x"fef42423",
x"2703a81d",
x"4789fec4",
x"00f70763",
x"fec42703",
x"18634791",
x"278300f7",
x"838dfe84",
x"fef42423",
x"2783a031",
x"8385fe84",
x"fef42423",
x"fec42783",
x"26230785",
x"2703fef4",
x"0793fe84",
x"e2e33fe0",
x"2223fce7",
x"2783fe04",
x"e793fe44",
x"22230017",
x"2783fef4",
x"078efec4",
x"27038be1",
x"8fd9fe44",
x"fef42223",
x"fe842783",
x"971317fd",
x"67c10067",
x"8ff917fd",
x"fe442703",
x"22238fd9",
x"77fdfef4",
x"50078793",
x"fe442703",
x"a011c398",
x"50b20001",
x"61455422",
x"11018082",
x"1000ce22",
x"fe042623",
x"e0000793",
x"07b74798",
x"8ff90002",
x"4785c781",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"d6067179",
x"1800d422",
x"fca42e23",
x"fe0407a3",
x"4703a821",
x"47a9fef4",
x"00f71463",
x"3d5d4535",
x"fef44783",
x"357d853e",
x"fdc42783",
x"00178713",
x"fce42e23",
x"0007c783",
x"fef407a3",
x"fef44783",
x"0001fbe9",
x"50b20001",
x"61455422",
x"11018082",
x"cc22ce06",
x"26231000",
x"2423fea4",
x"2583feb4",
x"2503fe84",
x"3545fec4",
x"40f20001",
x"61054462",
x"11018082",
x"cc22ce06",
x"26231000",
x"2503fea4",
x"3fbdfec4",
x"40f20001",
x"61054462",
x"11018082",
x"cc22ce06",
x"87aa1000",
x"fef407a3",
x"fef44783",
x"3d0d853e",
x"40f20001",
x"61054462",
x"71798082",
x"d422d606",
x"2e231800",
x"0513fca4",
x"3fc10300",
x"07800513",
x"262337e9",
x"a891fe04",
x"fdc42783",
x"242383f1",
x"2703fef4",
x"47a5fe84",
x"00e7cd63",
x"fe842783",
x"0ff7f793",
x"03078793",
x"0ff7f793",
x"3f71853e",
x"2783a819",
x"f793fe84",
x"87930ff7",
x"f7930377",
x"853e0ff7",
x"27833759",
x"0792fdc4",
x"fcf42e23",
x"fec42783",
x"26230785",
x"2703fef4",
x"479dfec4",
x"fae7d4e3",
x"00010001",
x"542250b2",
x"80826145",
x"d6067179",
x"1800d422",
x"fca42e23",
x"fe042623",
x"2783a815",
x"83f1fdc4",
x"fef42423",
x"fe842783",
x"0ff7f793",
x"03078793",
x"0ff7f793",
x"3735853e",
x"fdc42783",
x"2e230792",
x"2783fcf4",
x"0785fec4",
x"fef42623",
x"fec42703",
x"d4e3479d",
x"0001fce7",
x"50b20001",
x"61455422",
x"71798082",
x"d44ad622",
x"1800d24e",
x"fca42c23",
x"fcb42e23",
x"fe042623",
x"fdc42583",
x"0593e581",
x"a0110200",
x"24234581",
x"2503feb4",
x"2583fec4",
x"95aafe84",
x"feb42623",
x"fe842583",
x"c8631581",
x"25030005",
x"1eb3fd84",
x"4e0100b5",
x"2583a815",
x"d513fd84",
x"42fd0015",
x"fe842583",
x"40b285b3",
x"00b555b3",
x"fe842503",
x"fdc42283",
x"00a29eb3",
x"01d5eeb3",
x"fe842583",
x"fd842503",
x"00b51e33",
x"fdc42c23",
x"fdd42e23",
x"fdc42503",
x"746365c1",
x"45c100b5",
x"4581a011",
x"feb42423",
x"fec42503",
x"fe842583",
x"262395aa",
x"2583feb4",
x"1581fe84",
x"0005c863",
x"fd842503",
x"00b513b3",
x"a8154301",
x"fd842583",
x"0015d513",
x"25834e7d",
x"05b3fe84",
x"55b340be",
x"250300b5",
x"2e03fe84",
x"13b3fdc4",
x"e3b300ae",
x"25830075",
x"2503fe84",
x"1333fd84",
x"2c2300b5",
x"2e23fc64",
x"2503fc74",
x"05b7fdc4",
x"74630100",
x"45a100b5",
x"4581a011",
x"feb42423",
x"fec42503",
x"fe842583",
x"262395aa",
x"2583feb4",
x"1581fe84",
x"0005c863",
x"fd842503",
x"00b518b3",
x"a8154801",
x"fd842583",
x"0015d513",
x"2583437d",
x"05b3fe84",
x"55b340b3",
x"250300b5",
x"2303fe84",
x"18b3fdc4",
x"e8b300a3",
x"25830115",
x"2503fe84",
x"1833fd84",
x"2c2300b5",
x"2e23fd04",
x"2503fd14",
x"05b7fdc4",
x"74631000",
x"459100b5",
x"4581a011",
x"feb42423",
x"fec42503",
x"fe842583",
x"262395aa",
x"2583feb4",
x"1581fe84",
x"0005c863",
x"fd842503",
x"00b516b3",
x"a80d4601",
x"fd842583",
x"0015d513",
x"2583487d",
x"05b3fe84",
x"55b340b8",
x"250300b5",
x"2803fe84",
x"16b3fdc4",
x"8ecd00a8",
x"fe842583",
x"fd842503",
x"00b51633",
x"fcc42c23",
x"fcd42e23",
x"fdc42603",
x"400006b7",
x"00d67463",
x"a0114689",
x"24234681",
x"2603fed4",
x"2683fec4",
x"96b2fe84",
x"fed42623",
x"fe842683",
x"c8631681",
x"26030006",
x"17b3fd84",
x"470100d6",
x"2683a80d",
x"d613fd84",
x"45fd0016",
x"fe842683",
x"40d586b3",
x"00d656b3",
x"fe842603",
x"fdc42583",
x"00c597b3",
x"26838fd5",
x"2603fe84",
x"1733fd84",
x"2c2300d6",
x"2e23fce4",
x"2703fcf4",
x"2783fd84",
x"4f13fdc4",
x"cf93fff7",
x"d913fff7",
x"498101ff",
x"0ff97793",
x"2783873e",
x"97bafec4",
x"5432853e",
x"59925922",
x"80826145",
x"d7067171",
x"d326d522",
x"cf4ed14a",
x"cb56cd52",
x"c75ec95a",
x"c366c562",
x"deeec16a",
x"2c231900",
x"2e23f8a4",
x"2823f8b4",
x"2a23f8c4",
x"2623f8d4",
x"2703f8e4",
x"2783f944",
x"ee63f9c4",
x"270300e7",
x"2783f944",
x"1a63f9c4",
x"270302f7",
x"2783f904",
x"f463f984",
x"278302e7",
x"cb89f8c4",
x"f8c42683",
x"f9842703",
x"f9c42783",
x"c2dcc298",
x"48014781",
x"f8f42023",
x"f9042223",
x"2703a681",
x"2783f904",
x"e3f9f944",
x"f9042783",
x"f9442703",
x"e7958fd9",
x"fa0403a3",
x"fa744783",
x"0ff7f793",
x"87ba873e",
x"b7930785",
x"f7930037",
x"c3990ff7",
x"a01187ba",
x"f7934781",
x"03a30ff7",
x"2703faf4",
x"4785f904",
x"02f71763",
x"f9442783",
x"2783e39d",
x"c799f8c4",
x"f8c42783",
x"47014681",
x"c3d8c394",
x"f9842783",
x"f9c42803",
x"f8f42023",
x"f9042223",
x"2703a4f1",
x"2783f984",
x"eba9f9c4",
x"f8c42783",
x"2703c78d",
x"2783f984",
x"86baf9c4",
x"f9042703",
x"f9442783",
x"f7b387ba",
x"883e02f6",
x"27834881",
x"a023f8c4",
x"a2230107",
x"27030117",
x"2783f984",
x"86baf9c4",
x"f9042703",
x"f9442783",
x"d7b387ba",
x"202302f6",
x"2223f8f4",
x"ac8df804",
x"f9042503",
x"f9442583",
x"87aa390d",
x"0ff7f493",
x"f9842503",
x"f9c42583",
x"87aa310d",
x"0ff7f793",
x"40f487b3",
x"0ff7f793",
x"0fa30785",
x"4783faf4",
x"8713fbf4",
x"4863fe07",
x"27830007",
x"da33f9c4",
x"4a8100e7",
x"2703a01d",
x"1693f9c4",
x"477d0017",
x"97338f1d",
x"268300e6",
x"da33f984",
x"6a3300f6",
x"27030147",
x"5ab3f9c4",
x"282300f7",
x"2a23fb44",
x"4783fb54",
x"0713fbf4",
x"07b30400",
x"871340f7",
x"4863fe07",
x"27830007",
x"99b3f984",
x"490100e7",
x"2703a01d",
x"5693f984",
x"477d0017",
x"d7338f1d",
x"268300e6",
x"99b3f9c4",
x"69b300f6",
x"27030137",
x"1933f984",
x"2c2300f7",
x"2e23f924",
x"4781f934",
x"24234801",
x"2623faf4",
x"aa1dfb04",
x"fb042783",
x"270383fd",
x"1c93fb44",
x"ecb30017",
x"27830197",
x"9c13fb04",
x"27830017",
x"83fdf9c4",
x"f6f42c23",
x"f6042e23",
x"f7842683",
x"f7c42703",
x"67b387b6",
x"282300fc",
x"87bafaf4",
x"00fce7b3",
x"faf42a23",
x"f9842783",
x"270383fd",
x"1d93f9c4",
x"edb30017",
x"278301b7",
x"9d13f984",
x"27830017",
x"8b85fa84",
x"f6f42823",
x"fac42783",
x"2a238b81",
x"2683f6f4",
x"2703f704",
x"87b6f744",
x"00fd67b3",
x"f8f42c23",
x"e7b387ba",
x"2e2300fd",
x"2703f8f4",
x"2783f904",
x"2503f944",
x"2583fb04",
x"0633fb44",
x"883240a7",
x"01073833",
x"40b786b3",
x"410687b3",
x"557d86be",
x"073355fd",
x"883a00a6",
x"00c83833",
x"00b687b3",
x"00f806b3",
x"d69387b6",
x"242341f7",
x"87fdf6d4",
x"f6f42623",
x"f6842783",
x"f6c42803",
x"faf42423",
x"fb042623",
x"f9042703",
x"fa842783",
x"20238ff9",
x"2703f6f4",
x"2783f944",
x"8ff9fac4",
x"f6f42223",
x"fb042603",
x"fb442683",
x"f6042803",
x"f6442883",
x"073385c2",
x"85ba40b6",
x"00b635b3",
x"87b38546",
x"86b340a6",
x"87b640b7",
x"fae42823",
x"faf42a23",
x"fbf44783",
x"fff78713",
x"fae40fa3",
x"ec0790e3",
x"f8c42783",
x"2683cb89",
x"2703f8c4",
x"2783fb04",
x"c298fb44",
x"2783c2dc",
x"83fdf984",
x"f9c42703",
x"00171b93",
x"0177ebb3",
x"f9842783",
x"00179b13",
x"fa842783",
x"2c238b85",
x"2783f4f4",
x"8b81fac4",
x"f4f42e23",
x"f5842683",
x"f5c42703",
x"67b387b6",
x"202300fb",
x"87baf8f4",
x"00fbe7b3",
x"f8f42223",
x"f8042703",
x"f8442783",
x"85be853a",
x"542a50ba",
x"590a549a",
x"4a6a49fa",
x"4b4a4ada",
x"4c2a4bba",
x"4d0a4c9a",
x"614d5df6",
x"11018082",
x"cc22ce06",
x"24231000",
x"2623fea4",
x"2023feb4",
x"2223fec4",
x"4701fed4",
x"fe042603",
x"fe442683",
x"fe842503",
x"fec42583",
x"872a3ed5",
x"853a87ae",
x"40f285be",
x"61054462",
x"11018082",
x"1000ce22",
x"fea42623",
x"feb42423",
x"fe842783",
x"00079703",
x"fec42783",
x"00e79023",
x"fe842783",
x"00279703",
x"fec42783",
x"00e79123",
x"44720001",
x"80826105",
x"c686715d",
x"0880c4a2",
x"faa42e23",
x"fab42c23",
x"1b2387b2",
x"47d1faf4",
x"fef42223",
x"fbc42703",
x"fe442783",
x"02f757b3",
x"202317f9",
x"2703fef4",
x"2783fb84",
x"078efe04",
x"2e2397ba",
x"2783fcf4",
x"2423fdc4",
x"2703fcf4",
x"2783fc84",
x"078afe04",
x"2c2397ba",
x"2783fcf4",
x"2a23fb84",
x"2783fcf4",
x"a023fd44",
x"27030007",
x"2783fc84",
x"c3d8fd44",
x"fd442783",
x"912343dc",
x"27830007",
x"43dcfd44",
x"07137761",
x"90230807",
x"278300e7",
x"07a1fb84",
x"faf42c23",
x"fc842783",
x"24230791",
x"77e1fcf4",
x"fff7c793",
x"fcf41323",
x"122357fd",
x"0693fcf4",
x"0613fc84",
x"0593fb84",
x"2783fc44",
x"2703fd84",
x"2503fdc4",
x"2a91fd44",
x"fe042623",
x"2783a8ad",
x"9713fec4",
x"83410107",
x"fb645783",
x"07c28fb9",
x"8bbd83c1",
x"fcf41823",
x"fd045783",
x"9713078e",
x"83410107",
x"fec42783",
x"83c107c2",
x"07c28b9d",
x"8fd983c1",
x"fcf41723",
x"fce41783",
x"971307a2",
x"87410107",
x"fce41783",
x"07c28fd9",
x"122387c1",
x"0693fcf4",
x"0613fc84",
x"0593fb84",
x"2783fc44",
x"2703fd84",
x"2503fdc4",
x"20c5fd44",
x"fec42783",
x"26230785",
x"2703fef4",
x"2783fec4",
x"60e3fe04",
x"2783f8f7",
x"439cfd44",
x"fef42423",
x"26234785",
x"a841fef4",
x"fe042703",
x"57b34795",
x"270302f7",
x"7063fec4",
x"278302f7",
x"8713fec4",
x"26230017",
x"2703fee4",
x"4358fe84",
x"87c107c2",
x"00f71123",
x"2783a8a1",
x"8713fec4",
x"26230017",
x"9713fee4",
x"83410107",
x"fb645783",
x"19238fb9",
x"2783fcf4",
x"07c2fec4",
x"07a283c1",
x"83c107c2",
x"7007f793",
x"83c107c2",
x"fd245703",
x"07c28fd9",
x"969383c1",
x"86c10107",
x"fe842783",
x"671143dc",
x"8f75177d",
x"87410742",
x"00e79123",
x"fe842783",
x"2423439c",
x"2783fef4",
x"439cfe84",
x"4601f7b5",
x"5b400593",
x"fd442503",
x"f5bf60ef",
x"fca42a23",
x"fd442783",
x"40b6853e",
x"61614426",
x"71398082",
x"dc22de06",
x"2e230080",
x"2c23fca4",
x"2a23fcb4",
x"2823fcc4",
x"2623fcd4",
x"2423fce4",
x"2783fcf4",
x"439cfd44",
x"270307a1",
x"e463fcc4",
x"478100e7",
x"2783a895",
x"439cfd04",
x"27030791",
x"e463fc84",
x"478100e7",
x"2783a085",
x"439cfd44",
x"fef42623",
x"fd442783",
x"8713439c",
x"27830087",
x"c398fd44",
x"fdc42783",
x"27834398",
x"c398fec4",
x"fdc42783",
x"fec42703",
x"2783c398",
x"4398fd04",
x"fec42783",
x"2783c3d8",
x"439cfd04",
x"00478713",
x"fd042783",
x"2783c398",
x"43dcfec4",
x"fd842583",
x"3b01853e",
x"fec42783",
x"50f2853e",
x"61215462",
x"715d8082",
x"c4a2c686",
x"0880c2a6",
x"faa42e23",
x"fab42c23",
x"fe041623",
x"fe041523",
x"142357fd",
x"1323fef4",
x"1b23fe04",
x"4505fc04",
x"43b010ef",
x"971387aa",
x"87410107",
x"fbc42783",
x"00e79023",
x"10ef4509",
x"87aa4250",
x"01079713",
x"27838741",
x"9123fbc4",
x"450d00e7",
x"40f010ef",
x"971387aa",
x"87410107",
x"fbc42783",
x"00e79223",
x"10ef4511",
x"87aa3f90",
x"2783873e",
x"cfd8fbc4",
x"10ef4515",
x"87aa3e90",
x"2783873e",
x"d398fbc4",
x"fbc42783",
x"e789539c",
x"fbc42783",
x"d398471d",
x"fbc42783",
x"00079783",
x"2783eb8d",
x"9783fbc4",
x"e7850027",
x"fbc42783",
x"00479783",
x"2783ef99",
x"9023fbc4",
x"27830007",
x"9123fbc4",
x"27830007",
x"0713fbc4",
x"92230660",
x"278300e7",
x"9703fbc4",
x"47850007",
x"04f71063",
x"fbc42783",
x"00279783",
x"2783eb95",
x"9783fbc4",
x"e78d0047",
x"fbc42783",
x"0713670d",
x"90234157",
x"278300e7",
x"670dfbc4",
x"41570713",
x"00e79123",
x"fbc42783",
x"06600713",
x"00e79223",
x"fbc42783",
x"80000737",
x"12070713",
x"2783c798",
x"0713fbc4",
x"cf987d00",
x"fbc42783",
x"04079023",
x"fe041723",
x"5783a035",
x"4705fee4",
x"00f717b3",
x"2783873e",
x"539cfbc4",
x"c7918ff9",
x"fea45783",
x"15230785",
x"5783fef4",
x"0785fee4",
x"fef41723",
x"fee45703",
x"f8e34789",
x"1723fce7",
x"a081fe04",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"56834f90",
x"5703fea4",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fbc42783",
x"573397ba",
x"cf9802d6",
x"fee45783",
x"17230785",
x"5783fef4",
x"dfddfee4",
x"fe041723",
x"5783a071",
x"4705fee4",
x"00f717b3",
x"2783873e",
x"539cfbc4",
x"c7b58ff9",
x"fe042023",
x"2703a899",
x"87bafe04",
x"97ba0792",
x"873e078a",
x"fbc42783",
x"478c97ba",
x"fbc42783",
x"57834f98",
x"0633fec4",
x"270302f7",
x"87bafe04",
x"97ba0792",
x"873e078a",
x"fbc42783",
x"00e786b3",
x"fee45783",
x"87330785",
x"078a00c5",
x"c79897b6",
x"fe042783",
x"20230785",
x"2783fef4",
x"d7c5fe04",
x"fec45783",
x"16230785",
x"5783fef4",
x"0785fee4",
x"fef41723",
x"fee45703",
x"f8e34789",
x"1723f6e7",
x"aaa9fe04",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"8b85539c",
x"2783cbb1",
x"4f94fbc4",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"570347cc",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fbc42783",
x"960397ba",
x"57030007",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fbc42783",
x"00e784b3",
x"34bd8536",
x"d0dc87aa",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"8b89539c",
x"2783cbb5",
x"4f88fbc4",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"57034b8c",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fbc42783",
x"978397ba",
x"86be0007",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"00279783",
x"e63307c2",
x"570300f6",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fbc42783",
x"879397ba",
x"86be0287",
x"838f70ef",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"8b91539c",
x"2783cf9d",
x"4f94fbc4",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"00079583",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"863e4bdc",
x"10ef8536",
x"57834160",
x"0785fee4",
x"fef41723",
x"fee45783",
x"ea0782e3",
x"fbc42783",
x"e3d14fdc",
x"fc042e23",
x"fbc42783",
x"cfd84705",
x"2783a081",
x"4fd8fbc4",
x"078a87ba",
x"078697ba",
x"2783873e",
x"cfd8fbc4",
x"132010ef",
x"fbc42503",
x"ec1f60ef",
x"14a010ef",
x"16a010ef",
x"87ae872a",
x"fb842603",
x"85be853a",
x"19e010ef",
x"fca42e23",
x"fdc42783",
x"2783dfdd",
x"2c23fdc4",
x"2783fcf4",
x"e781fd84",
x"2c234785",
x"2783fcf4",
x"4fd8fbc4",
x"278346a9",
x"d7b3fd84",
x"078502f6",
x"02f70733",
x"fbc42783",
x"10efcfd8",
x"25030d40",
x"60effbc4",
x"10efe63f",
x"10ef0ec0",
x"242310c0",
x"2623fca4",
x"2783fcb4",
x"9783fbc4",
x"57030007",
x"85bafd64",
x"70ef853e",
x"87aac30f",
x"fcf41b23",
x"fbc42783",
x"00279783",
x"fd645703",
x"853e85ba",
x"c16f70ef",
x"1b2387aa",
x"2783fcf4",
x"9783fbc4",
x"57030047",
x"85bafd64",
x"70ef853e",
x"87aabfcf",
x"fcf41b23",
x"fbc42783",
x"07c24f9c",
x"570387c1",
x"85bafd64",
x"70ef853e",
x"87aabe0f",
x"fcf41b23",
x"fd645783",
x"0713673d",
x"81639f57",
x"673d06e7",
x"9f570713",
x"06f74463",
x"07136725",
x"8c63a027",
x"672502e7",
x"a0270713",
x"04f74a63",
x"07136721",
x"8563b057",
x"672102e7",
x"b0570713",
x"04f74063",
x"07136709",
x"87638f27",
x"671502e7",
x"eaf70713",
x"00e78a63",
x"1423a025",
x"a02dfe04",
x"14234785",
x"a00dfef4",
x"14234789",
x"a829fef4",
x"1423478d",
x"a809fef4",
x"14234791",
x"a029fef4",
x"132357fd",
x"0001fef4",
x"fe841783",
x"1c07c263",
x"fe041723",
x"5703a275",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fbc42783",
x"902397ba",
x"57030407",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fbc42783",
x"539c97ba",
x"cfb18b85",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"03a7d703",
x"fe841783",
x"800006b7",
x"00068693",
x"97b60786",
x"0007d783",
x"02f70763",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"04079703",
x"83410742",
x"07420705",
x"07428341",
x"90238741",
x"570304e7",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fbc42783",
x"539c97ba",
x"cfb18b89",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"03c7d703",
x"fe841783",
x"800006b7",
x"00c68693",
x"97b60786",
x"0007d783",
x"02f70763",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"04079703",
x"83410742",
x"07420705",
x"07428341",
x"90238741",
x"570304e7",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fbc42783",
x"539c97ba",
x"cfb18b91",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"03e7d703",
x"fe841783",
x"800006b7",
x"01868693",
x"97b60786",
x"0007d783",
x"02f70763",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"04079703",
x"83410742",
x"07420705",
x"07428341",
x"90238741",
x"570304e7",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fbc42783",
x"978397ba",
x"97130407",
x"83410107",
x"fe645783",
x"07c297ba",
x"132383c1",
x"5783fef4",
x"0785fee4",
x"fef41723",
x"fee45703",
x"800007b7",
x"0707a783",
x"e4f765e3",
x"5ba010ef",
x"873e87aa",
x"fe645783",
x"07c297ba",
x"132383c1",
x"2783fef4",
x"4f9cfbc4",
x"67a185be",
x"16078513",
x"276020ef",
x"fc842703",
x"fcc42783",
x"3e800613",
x"853a4681",
x"f0ef85be",
x"872ad6cf",
x"87ba87ae",
x"67a185be",
x"17878513",
x"24e020ef",
x"fb842603",
x"fc842503",
x"fcc42583",
x"633000ef",
x"85be87aa",
x"851367a1",
x"20ef1947",
x"26032300",
x"2503fb84",
x"2583fc84",
x"00effcc4",
x"87aa6150",
x"2783cb9d",
x"4fd8fbc4",
x"800007b7",
x"0707a783",
x"02f704b3",
x"fb842603",
x"fc842503",
x"fcc42583",
x"5ef000ef",
x"d7b387aa",
x"85be02f4",
x"851367a1",
x"20ef1ac7",
x"26031e80",
x"2503fb84",
x"2583fc84",
x"00effcc4",
x"872a5cd0",
x"e06347a5",
x"67a102e7",
x"1c478513",
x"1c6020ef",
x"fe641783",
x"83c107c2",
x"07c20785",
x"132383c1",
x"2783fef4",
x"4fd8fbc4",
x"800007b7",
x"0707a783",
x"02f707b3",
x"67a185be",
x"20478513",
x"196020ef",
x"859367a1",
x"67a121c7",
x"22878513",
x"186020ef",
x"859367a1",
x"67a12407",
x"25c78513",
x"176020ef",
x"859367a1",
x"67a12747",
x"27c78513",
x"166020ef",
x"fd645783",
x"67a185be",
x"29478513",
x"156020ef",
x"fbc42783",
x"8b85539c",
x"1723c7b1",
x"a81dfe04",
x"fee45683",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"03a7d783",
x"85b6863e",
x"851367a1",
x"20ef2b07",
x"578311c0",
x"0785fee4",
x"fef41723",
x"fee45703",
x"800007b7",
x"0707a783",
x"fcf760e3",
x"fbc42783",
x"8b89539c",
x"1723c7b1",
x"a81dfe04",
x"fee45683",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"03c7d783",
x"85b6863e",
x"851367a1",
x"20ef2cc7",
x"57830c80",
x"0785fee4",
x"fef41723",
x"fee45703",
x"800007b7",
x"0707a783",
x"fcf760e3",
x"fbc42783",
x"8b91539c",
x"1723c7b1",
x"a81dfe04",
x"fee45683",
x"fee45703",
x"079287ba",
x"078a97ba",
x"2783873e",
x"97bafbc4",
x"03e7d783",
x"85b6863e",
x"851367a1",
x"20ef2e87",
x"57830740",
x"0785fee4",
x"fef41723",
x"fee45703",
x"800007b7",
x"0707a783",
x"fcf760e3",
x"fe041723",
x"5683a81d",
x"5703fee4",
x"87bafee4",
x"97ba0792",
x"873e078a",
x"fbc42783",
x"d78397ba",
x"863e0387",
x"67a185b6",
x"30478513",
x"02a020ef",
x"fee45783",
x"17230785",
x"5703fef4",
x"07b7fee4",
x"a7838000",
x"60e30707",
x"1783fcf7",
x"e791fe64",
x"851367a1",
x"20ef3207",
x"17830000",
x"5763fe64",
x"67a100f0",
x"36c78513",
x"7ef010ef",
x"fe641783",
x"0007d763",
x"851367a1",
x"10ef3807",
x"47817dd0",
x"40b6853e",
x"44964426",
x"80826161",
x"de067139",
x"0080dc22",
x"fca42e23",
x"fcb42c23",
x"fcc42a23",
x"fcd42823",
x"172387ba",
x"1723fcf4",
x"5783fe04",
x"873efce4",
x"8fd977fd",
x"fef41623",
x"fce41783",
x"2583863e",
x"2503fd44",
x"2469fdc4",
x"fce41783",
x"260386be",
x"2583fd44",
x"2503fd84",
x"2ae1fdc4",
x"fec41783",
x"2583863e",
x"2503fd84",
x"20edfdc4",
x"873e87aa",
x"fee45783",
x"853a85be",
x"e4bf60ef",
x"172387aa",
x"2683fef4",
x"2603fd04",
x"2583fd44",
x"2503fd84",
x"24e5fdc4",
x"fec41783",
x"2583863e",
x"2503fd84",
x"284dfdc4",
x"873e87aa",
x"fee45783",
x"853a85be",
x"e13f60ef",
x"172387aa",
x"2683fef4",
x"2603fd04",
x"2583fd44",
x"2503fd84",
x"26adfdc4",
x"fec41783",
x"2583863e",
x"2503fd84",
x"28adfdc4",
x"873e87aa",
x"fee45783",
x"853a85be",
x"ddbf60ef",
x"172387aa",
x"2683fef4",
x"2603fd04",
x"2583fd44",
x"2503fd84",
x"2181fdc4",
x"fec41783",
x"2583863e",
x"2503fd84",
x"2089fdc4",
x"873e87aa",
x"fee45783",
x"853a85be",
x"da3f60ef",
x"172387aa",
x"5783fef4",
x"07b3fce4",
x"07c240f0",
x"07c283c1",
x"863e87c1",
x"fd442583",
x"fdc42503",
x"17832271",
x"853efee4",
x"546250f2",
x"80826121",
x"de227139",
x"26230080",
x"2423fca4",
x"87b2fcb4",
x"fcf41323",
x"fe042623",
x"fe042423",
x"fc042c23",
x"fe041323",
x"fe042023",
x"2e23a879",
x"a049fc04",
x"fe042703",
x"fcc42783",
x"02f70733",
x"fdc42783",
x"078a97ba",
x"fc842703",
x"439c97ba",
x"fcf42c23",
x"fec42703",
x"fd842783",
x"262397ba",
x"1783fef4",
x"2703fc64",
x"dc63fec4",
x"578300e7",
x"07a9fe64",
x"83c107c2",
x"fef41323",
x"fe042623",
x"2703a00d",
x"2783fd84",
x"a7b3fe84",
x"f79300e7",
x"873e0ff7",
x"fe645783",
x"07c297ba",
x"132383c1",
x"2783fef4",
x"2423fd84",
x"2783fef4",
x"0785fdc4",
x"fcf42e23",
x"fdc42703",
x"fcc42783",
x"f6f76ce3",
x"fe042783",
x"20230785",
x"2703fef4",
x"2783fe04",
x"6ee3fcc4",
x"1783f4f7",
x"853efe64",
x"61215472",
x"71798082",
x"1800d622",
x"fca42e23",
x"fcb42c23",
x"fcc42a23",
x"192387b6",
x"2623fcf4",
x"a0b5fe04",
x"fe042423",
x"2703a881",
x"2783fec4",
x"0733fdc4",
x"278302f7",
x"97bafe84",
x"27030786",
x"97bafd44",
x"00079783",
x"1703863e",
x"2683fd24",
x"2783fec4",
x"86b3fdc4",
x"278302f6",
x"97b6fe84",
x"2683078a",
x"97b6fd84",
x"02e60733",
x"2783c398",
x"0785fe84",
x"fef42423",
x"fe842703",
x"fdc42783",
x"faf765e3",
x"fec42783",
x"26230785",
x"2703fef4",
x"2783fec4",
x"67e3fdc4",
x"0001f8f7",
x"54320001",
x"80826145",
x"d6227179",
x"2e231800",
x"2c23fca4",
x"87b2fcb4",
x"fcf41b23",
x"fe042623",
x"2423a8b5",
x"a085fe04",
x"fec42703",
x"fdc42783",
x"02f70733",
x"fe842783",
x"078697ba",
x"fd842703",
x"978397ba",
x"97130007",
x"83410107",
x"fd645783",
x"969397ba",
x"82c10107",
x"fec42703",
x"fdc42783",
x"02f70733",
x"fe842783",
x"078697ba",
x"fd842703",
x"971397ba",
x"87410106",
x"00e79023",
x"fe842783",
x"24230785",
x"2703fef4",
x"2783fe84",
x"6de3fdc4",
x"2783f8f7",
x"0785fec4",
x"fef42623",
x"fec42703",
x"fdc42783",
x"f6f76fe3",
x"00010001",
x"61455432",
x"71798082",
x"1800d622",
x"fca42e23",
x"fcb42c23",
x"fcc42a23",
x"fcd42823",
x"fe042623",
x"2783a069",
x"078afec4",
x"fd842703",
x"a02397ba",
x"24230007",
x"a8b9fe04",
x"fec42783",
x"2703078a",
x"97bafd84",
x"27034394",
x"2783fec4",
x"0733fdc4",
x"278302f7",
x"97bafe84",
x"27030786",
x"97bafd44",
x"00079783",
x"2783863e",
x"0786fe84",
x"fd042703",
x"978397ba",
x"07330007",
x"278302f6",
x"078afec4",
x"fd842603",
x"973697b2",
x"2783c398",
x"0785fe84",
x"fef42423",
x"fe842703",
x"fdc42783",
x"f8f76ee3",
x"fec42783",
x"26230785",
x"2703fef4",
x"2783fec4",
x"68e3fdc4",
x"0001f6f7",
x"54320001",
x"80826145",
x"d6227179",
x"2e231800",
x"2c23fca4",
x"2a23fcb4",
x"2823fcc4",
x"2623fcd4",
x"a8f9fe04",
x"fe042423",
x"2703a0c9",
x"2783fec4",
x"0733fdc4",
x"278302f7",
x"97bafe84",
x"2703078a",
x"97bafd84",
x"0007a023",
x"fe042223",
x"2703a061",
x"2783fec4",
x"0733fdc4",
x"278302f7",
x"97bafe84",
x"2703078a",
x"97bafd84",
x"27034394",
x"2783fec4",
x"0733fdc4",
x"278302f7",
x"97bafe44",
x"27030786",
x"97bafd44",
x"00079783",
x"2703863e",
x"2783fe44",
x"0733fdc4",
x"278302f7",
x"97bafe84",
x"27030786",
x"97bafd04",
x"00079783",
x"02f60733",
x"fec42603",
x"fdc42783",
x"02f60633",
x"fe842783",
x"078a97b2",
x"fd842603",
x"973697b2",
x"2783c398",
x"0785fe44",
x"fef42223",
x"fe442703",
x"fdc42783",
x"f6f769e3",
x"fe842783",
x"24230785",
x"2703fef4",
x"2783fe84",
x"6ce3fdc4",
x"2783f2f7",
x"0785fec4",
x"fef42623",
x"fec42703",
x"fdc42783",
x"f0f76ee3",
x"00010001",
x"61455432",
x"71798082",
x"1800d622",
x"fca42e23",
x"fcb42c23",
x"fcc42a23",
x"fcd42823",
x"fe042623",
x"2423a8fd",
x"a0cdfe04",
x"fec42703",
x"fdc42783",
x"02f70733",
x"fe842783",
x"078a97ba",
x"fd842703",
x"a02397ba",
x"22230007",
x"a065fe04",
x"fec42703",
x"fdc42783",
x"02f70733",
x"fe442783",
x"078697ba",
x"fd442703",
x"978397ba",
x"86be0007",
x"fe442703",
x"fdc42783",
x"02f70733",
x"fe842783",
x"078697ba",
x"fd042703",
x"978397ba",
x"87b30007",
x"202302f6",
x"2703fef4",
x"2783fec4",
x"0733fdc4",
x"278302f7",
x"97bafe84",
x"2703078a",
x"97bafd84",
x"86be439c",
x"fe042783",
x"f7138789",
x"278300f7",
x"8795fe04",
x"07f7f793",
x"02f707b3",
x"270396be",
x"2783fec4",
x"0733fdc4",
x"278302f7",
x"97bafe84",
x"2703078a",
x"97bafd84",
x"c3988736",
x"fe442783",
x"22230785",
x"2703fef4",
x"2783fe44",
x"69e3fdc4",
x"2783f4f7",
x"0785fe84",
x"fef42423",
x"fe842703",
x"fdc42783",
x"f0f76ce3",
x"fec42783",
x"26230785",
x"2703fef4",
x"2783fec4",
x"6ee3fdc4",
x"0001eef7",
x"54320001",
x"80826145",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"00013047",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"32079073",
x"44720001",
x"80826105",
x"ce221101",
x"27f31000",
x"2623b000",
x"2783fef4",
x"863efec4",
x"87324681",
x"853a87b6",
x"447285be",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"0001b007",
x"61054472",
x"11018082",
x"1000ce22",
x"b02027f3",
x"fef42623",
x"fec42783",
x"4681863e",
x"87b68732",
x"85be853a",
x"61054472",
x"11018082",
x"1000ce22",
x"b03027f3",
x"fef42623",
x"fec42783",
x"4681863e",
x"87b68732",
x"85be853a",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"b0379073",
x"44720001",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"00013237",
x"61054472",
x"11018082",
x"1000ce22",
x"c00027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce221101",
x"27f31000",
x"2623c800",
x"2783fef4",
x"853efec4",
x"61054472",
x"11018082",
x"1000ce22",
x"b04027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"0001b047",
x"61054472",
x"11018082",
x"1000ce22",
x"b05027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"0001b057",
x"61054472",
x"11018082",
x"1000ce22",
x"b06027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"0001b067",
x"61054472",
x"11018082",
x"1000ce22",
x"b07027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"0001b077",
x"61054472",
x"11018082",
x"1000ce22",
x"b08027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"0001b087",
x"61054472",
x"11018082",
x"1000ce22",
x"b09027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"0001b097",
x"61054472",
x"11018082",
x"1000ce22",
x"b0a027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"0001b0a7",
x"61054472",
x"11018082",
x"1000ce22",
x"b0b027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"0001b0b7",
x"61054472",
x"11018082",
x"1000ce22",
x"b0c027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"0001b0c7",
x"61054472",
x"11018082",
x"1000ce22",
x"b0d027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"0001b0d7",
x"61054472",
x"11018082",
x"1000ce22",
x"b0e027f3",
x"fef42623",
x"fec42783",
x"4472853e",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"0001b0e7",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"32479073",
x"44720001",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"00013257",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"32679073",
x"44720001",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"00013277",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"32879073",
x"44720001",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"00013297",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"32a79073",
x"44720001",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"000132b7",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"32c79073",
x"44720001",
x"80826105",
x"ce221101",
x"26231000",
x"2783fea4",
x"9073fec4",
x"000132d7",
x"61054472",
x"11018082",
x"1000ce22",
x"fea42623",
x"fec42783",
x"32e79073",
x"44720001",
x"80826105",
x"d6067179",
x"1800d422",
x"26233151",
x"3195fea4",
x"fea42423",
x"222339a5",
x"2703fea4",
x"2783fec4",
x"0363fe44",
x"b7cd00f7",
x"27830001",
x"2c23fe84",
x"2783fcf4",
x"2e23fe44",
x"2703fcf4",
x"2783fd84",
x"853afdc4",
x"50b285be",
x"61455422",
x"11418082",
x"c422c606",
x"376d0800",
x"87ae872a",
x"82e1a423",
x"82f1a623",
x"3e254501",
x"40b20001",
x"01414422",
x"11418082",
x"c422c606",
x"557d0800",
x"3749360d",
x"87ae872a",
x"82e1a823",
x"82f1aa23",
x"40b20001",
x"01414422",
x"11018082",
x"1000ce22",
x"8301a603",
x"8341a683",
x"8281a503",
x"82c1a583",
x"40a60733",
x"3833883a",
x"87b30106",
x"86b340b6",
x"87b64107",
x"fee42423",
x"fef42623",
x"fe842703",
x"fec42783",
x"85be853a",
x"61054472",
x"71798082",
x"d422d606",
x"2c231800",
x"2e23fca4",
x"2a23fcb4",
x"2683fcc4",
x"8736fd44",
x"863a4781",
x"250386be",
x"2583fd84",
x"e0effdc4",
x"872aef0f",
x"262387ae",
x"2783fee4",
x"853efec4",
x"542250b2",
x"80826145",
x"ce061101",
x"1000cc22",
x"fea42623",
x"feb42423",
x"3c994501",
x"34b5557d",
x"345d4501",
x"36114501",
x"3e294521",
x"3ebd4501",
x"3b714541",
x"366d4501",
x"02000513",
x"45013375",
x"05133ed1",
x"3b750400",
x"3efd4501",
x"08000513",
x"450133f1",
x"05133125",
x"3bf11000",
x"39894501",
x"20000513",
x"450133f5",
x"051339b5",
x"3bf54000",
x"315d4501",
x"85136785",
x"35298007",
x"31f94501",
x"3d316505",
x"39ed4501",
x"353d6509",
x"331d4501",
x"35816511",
x"fe842503",
x"f8dfd0ef",
x"d0ef4529",
x"4529ee1f",
x"f81fd0ef",
x"d0ef4529",
x"2783ed5f",
x"4705fec4",
x"00e78023",
x"40f20001",
x"61054462",
x"11018082",
x"cc22ce06",
x"26231000",
x"2783fea4",
x"8023fec4",
x"67a10007",
x"3e478513",
x"e87fd0ef",
x"872a32d1",
x"87ba87ae",
x"d0ef853e",
x"4529eb5f",
x"e8ffd0ef",
x"872a32fd",
x"87ba87ae",
x"d0ef853e",
x"4529ea1f",
x"e7bfd0ef",
x"872a3afd",
x"87ba87ae",
x"d0ef853e",
x"4529e8df",
x"e67fd0ef",
x"87aa3c9d",
x"d0ef853e",
x"4529e7df",
x"e57fd0ef",
x"87aa3c69",
x"d0ef853e",
x"4529e6df",
x"e47fd0ef",
x"87aa3c7d",
x"d0ef853e",
x"4529e5df",
x"e37fd0ef",
x"87aa34cd",
x"d0ef853e",
x"4529e4df",
x"e27fd0ef",
x"87aa3619",
x"d0ef853e",
x"4529e3df",
x"e17fd0ef",
x"87aa362d",
x"d0ef853e",
x"4529e2df",
x"e07fd0ef",
x"87aa36b9",
x"d0ef853e",
x"4529e1df",
x"df7fd0ef",
x"87aa3e8d",
x"d0ef853e",
x"4529e0df",
x"de7fd0ef",
x"87aa3e59",
x"d0ef853e",
x"4529dfdf",
x"dd7fd0ef",
x"87aa3e6d",
x"d0ef853e",
x"4529dedf",
x"dc7fd0ef",
x"87aa3ef9",
x"d0ef853e",
x"4529dddf",
x"db7fd0ef",
x"d0ef4529",
x"0001db1f",
x"446240f2",
x"80826105",
x"d6227179",
x"2e231800",
x"87aefca4",
x"fcc42a23",
x"fcf41d23",
x"fe042623",
x"fe042423",
x"fe042023",
x"fdc42783",
x"2e2317fd",
x"2423fcf4",
x"a285fe04",
x"fe842783",
x"2223c7a5",
x"a03dfe04",
x"fe042703",
x"fe442783",
x"2683973e",
x"2783fec4",
x"97b6fe44",
x"fd442683",
x"470397b6",
x"80230007",
x"278300e7",
x"0785fe44",
x"fef42223",
x"fe442703",
x"fe842783",
x"fcf766e3",
x"fec42703",
x"fe442783",
x"270397ba",
x"97bafd44",
x"02c00713",
x"00e78023",
x"fe842703",
x"fec42783",
x"078597ba",
x"fef42623",
x"fda41783",
x"83c107c2",
x"07c20785",
x"1d2383c1",
x"5783fcf4",
x"8b9dfda4",
x"8663471d",
x"471d0ae7",
x"0cf74863",
x"45634719",
x"47150cf7",
x"06e7d863",
x"45634709",
x"d96300f7",
x"a85d0007",
x"ffd78713",
x"e7634785",
x"a0350ae7",
x"fda41783",
x"07c2878d",
x"07c287c1",
x"8b8d83c1",
x"80000737",
x"02470713",
x"97ba078a",
x"2023439c",
x"4791fef4",
x"fef42423",
x"1783a049",
x"878dfda4",
x"87c107c2",
x"83c107c2",
x"07378b8d",
x"07138000",
x"078a0347",
x"439c97ba",
x"fef42023",
x"242347a1",
x"a8a1fef4",
x"fda41783",
x"07c2878d",
x"07c287c1",
x"8b8d83c1",
x"80000737",
x"04470713",
x"97ba078a",
x"2023439c",
x"47a1fef4",
x"fef42423",
x"1783a03d",
x"878dfda4",
x"87c107c2",
x"83c107c2",
x"07378b8d",
x"07138000",
x"078a0547",
x"439c97ba",
x"fef42023",
x"242347a1",
x"a011fef4",
x"27030001",
x"2783fec4",
x"97bafe84",
x"27030785",
x"e9e3fdc4",
x"2783e8e7",
x"0785fdc4",
x"fcf42e23",
x"2703a829",
x"2783fd44",
x"97bafec4",
x"00078023",
x"fec42783",
x"26230785",
x"2703fef4",
x"2783fec4",
x"60e3fdc4",
x"0001fef7",
x"54320001",
x"80826145",
x"d6227179",
x"87aa1800",
x"fcf40fa3",
x"fdf44783",
x"0307b793",
x"0017b793",
x"0ff7f713",
x"fdf44783",
x"03a7b793",
x"0ff7f793",
x"f7938ff9",
x"07a30ff7",
x"4783fef4",
x"853efef4",
x"61455432",
x"71798082",
x"d422d606",
x"2e231800",
x"2c23fca4",
x"2783fcb4",
x"439cfdc4",
x"fef42623",
x"fe042423",
x"2783ac3d",
x"c783fec4",
x"03a30007",
x"4703fef4",
x"0793fe74",
x"186302c0",
x"278300f7",
x"0785fec4",
x"fef42623",
x"2703a43d",
x"479dfe84",
x"1ee7ed63",
x"fe842783",
x"00279713",
x"879367a1",
x"97ba4d07",
x"8782439c",
x"fe744783",
x"3fa9853e",
x"c78987aa",
x"24234791",
x"a0a1fef4",
x"fe744703",
x"02b00793",
x"00f70863",
x"fe744703",
x"02d00793",
x"00f71663",
x"24234789",
x"a025fef4",
x"fe744703",
x"02e00793",
x"00f71663",
x"24234795",
x"a811fef4",
x"24234785",
x"2783fef4",
x"0791fd84",
x"07054398",
x"2783c398",
x"439cfd84",
x"00178713",
x"fd842783",
x"a259c398",
x"fe744783",
x"35fd853e",
x"cb9987aa",
x"24234791",
x"2783fef4",
x"07a1fd84",
x"07054398",
x"a29dc398",
x"fe744703",
x"02e00793",
x"00f71c63",
x"24234795",
x"2783fef4",
x"07a1fd84",
x"07054398",
x"a299c398",
x"24234785",
x"2783fef4",
x"07a1fd84",
x"07054398",
x"aa0dc398",
x"fe744703",
x"02e00793",
x"00f71c63",
x"24234795",
x"2783fef4",
x"07c1fd84",
x"07054398",
x"a221c398",
x"fe744783",
x"3dad853e",
x"9e6387aa",
x"47850e07",
x"fef42423",
x"fd842783",
x"439807c1",
x"c3980705",
x"4703a0dd",
x"0793fe74",
x"08630450",
x"470300f7",
x"0793fe74",
x"1c630650",
x"478d00f7",
x"fef42423",
x"fd842783",
x"439807d1",
x"c3980705",
x"4783a87d",
x"853efe74",
x"87aa3535",
x"4785ebcd",
x"fef42423",
x"fd842783",
x"439807d1",
x"c3980705",
x"4703a879",
x"0793fe74",
x"086302b0",
x"470300f7",
x"0793fe74",
x"1c6302d0",
x"479900f7",
x"fef42423",
x"fd842783",
x"439807b1",
x"c3980705",
x"4785a8a5",
x"fef42423",
x"fd842783",
x"439807b1",
x"c3980705",
x"4783a095",
x"853efe74",
x"87aa33f1",
x"479dcb99",
x"fef42423",
x"fd842783",
x"439807e1",
x"c3980705",
x"4785a091",
x"fef42423",
x"fd842783",
x"439807e1",
x"c3980705",
x"4783a805",
x"853efe74",
x"87aa3b61",
x"4785e38d",
x"fef42423",
x"fd842783",
x"43980791",
x"c3980705",
x"0001a039",
x"0001a031",
x"0001a021",
x"0001a011",
x"fec42783",
x"26230785",
x"2783fef4",
x"c783fec4",
x"c7910007",
x"fe842703",
x"1ae34785",
x"2783daf7",
x"2703fdc4",
x"c398fec4",
x"fe842783",
x"50b2853e",
x"61455422",
x"71798082",
x"1800d622",
x"fca42e23",
x"fdc42703",
x"e9634795",
x"278304e7",
x"9713fdc4",
x"67a10027",
x"4f078793",
x"439c97ba",
x"a7838782",
x"26238181",
x"a825fef4",
x"81c1a783",
x"fef42623",
x"07b7a03d",
x"a7838000",
x"26230687",
x"a005fef4",
x"800007b7",
x"06c7a783",
x"fef42623",
x"a783a809",
x"26238201",
x"a021fef4",
x"fe042623",
x"27830001",
x"853efec4",
x"61455432",
x"11018082",
x"cc22ce06",
x"07a31000",
x"4783fe04",
x"c791fef4",
x"851367a1",
x"00ef5087",
x"47834c90",
x"853efef4",
x"446240f2",
x"80826105",
x"d6227179",
x"2e231800",
x"2c23fca4",
x"2783fcb4",
x"2623fdc4",
x"a031fef4",
x"fec42783",
x"26230785",
x"2783fef4",
x"c783fec4",
x"cb810007",
x"fd842783",
x"fff78713",
x"fce42c23",
x"2703f3e5",
x"2783fec4",
x"07b3fdc4",
x"853e40f7",
x"61455432",
x"71798082",
x"1800d622",
x"fca42e23",
x"fe042623",
x"2703a03d",
x"87bafec4",
x"97ba078a",
x"863e0786",
x"fdc42783",
x"8693439c",
x"27030017",
x"c314fdc4",
x"0007c783",
x"879397b2",
x"2623fd07",
x"2783fef4",
x"439cfdc4",
x"0007c703",
x"02f00793",
x"00e7fb63",
x"fdc42783",
x"c703439c",
x"07930007",
x"fae30390",
x"2783fae7",
x"853efec4",
x"61455432",
x"71198082",
x"0100dea2",
x"f8a42e23",
x"f8b42c23",
x"f8c42a23",
x"f8d42823",
x"f8e42623",
x"f8f42423",
x"80c1a783",
x"fef42423",
x"f8842783",
x"0407f793",
x"a783c789",
x"24238101",
x"2783fef4",
x"8bc1f884",
x"2783c791",
x"9bf9f884",
x"f8f42423",
x"f9442703",
x"d8634785",
x"270300e7",
x"0793f944",
x"d4630240",
x"478100e7",
x"2783ac59",
x"8b85f884",
x"0793c781",
x"a0190300",
x"02000793",
x"fef401a3",
x"fe0407a3",
x"f8842783",
x"c3a58b89",
x"f9842783",
x"0207d263",
x"02d00793",
x"fef407a3",
x"f9842783",
x"40f007b3",
x"f8f42c23",
x"f9042783",
x"282317fd",
x"a825f8f4",
x"f8842783",
x"cb998b91",
x"02b00793",
x"fef407a3",
x"f9042783",
x"282317fd",
x"a831f8f4",
x"f8842783",
x"cb918ba1",
x"02000793",
x"fef407a3",
x"f9042783",
x"282317fd",
x"2783f8f4",
x"f793f884",
x"c7950207",
x"f9442703",
x"186347c1",
x"278300f7",
x"17f9f904",
x"f8f42823",
x"2703a819",
x"47a1f944",
x"00f71763",
x"f9042783",
x"282317fd",
x"2223f8f4",
x"2783fe04",
x"ebb9f984",
x"fe442783",
x"00178713",
x"fee42223",
x"97a217c1",
x"03000713",
x"fae78823",
x"2703a089",
x"2783f984",
x"77b3f944",
x"270302f7",
x"973efe84",
x"fe442783",
x"00178693",
x"fed42223",
x"00074703",
x"97a217c1",
x"fae78823",
x"f9842703",
x"f9442783",
x"02f757b3",
x"f8f42c23",
x"f9842783",
x"2703f3e9",
x"2783fe44",
x"d663f8c4",
x"278300e7",
x"2623fe44",
x"2703f8f4",
x"2783f904",
x"07b3f8c4",
x"282340f7",
x"2783f8f4",
x"8bc5f884",
x"a819e785",
x"f9c42783",
x"00178713",
x"f8e42e23",
x"02000713",
x"00e78023",
x"f9042783",
x"fff78713",
x"f8e42823",
x"fef040e3",
x"fef44783",
x"2783cb99",
x"8713f9c4",
x"2e230017",
x"4703f8e4",
x"8023fef4",
x"278300e7",
x"f793f884",
x"cfa10207",
x"f9442703",
x"1d6347a1",
x"278300f7",
x"8713f9c4",
x"2e230017",
x"0713f8e4",
x"80230300",
x"a82500e7",
x"f9442703",
x"186347c1",
x"278302f7",
x"8713f9c4",
x"2e230017",
x"0713f8e4",
x"80230300",
x"a70300e7",
x"278380c1",
x"8693f9c4",
x"2e230017",
x"4703f8d4",
x"80230217",
x"278300e7",
x"8bc1f884",
x"a819ef9d",
x"f9c42783",
x"00178713",
x"f8e42e23",
x"fe344703",
x"00e78023",
x"f9042783",
x"fff78713",
x"f8e42823",
x"fef040e3",
x"2783a819",
x"8713f9c4",
x"2e230017",
x"0713f8e4",
x"80230300",
x"278300e7",
x"8713f8c4",
x"2623fff7",
x"2703f8e4",
x"4ee3fe44",
x"a839fcf7",
x"f9c42783",
x"00178713",
x"f8e42e23",
x"fe442703",
x"97221741",
x"fb074703",
x"00e78023",
x"fe442783",
x"fff78713",
x"fee42223",
x"fcf04ce3",
x"2783a819",
x"8713f9c4",
x"2e230017",
x"0713f8e4",
x"80230200",
x"278300e7",
x"8713f904",
x"2823fff7",
x"40e3f8e4",
x"2783fef0",
x"853ef9c4",
x"61095476",
x"711d8082",
x"1080cea2",
x"faa42e23",
x"fab42c23",
x"fac42a23",
x"fad42823",
x"fae42623",
x"80c1a783",
x"fef42623",
x"fac42783",
x"0407f793",
x"a783c789",
x"26238101",
x"2223fef4",
x"2423fe04",
x"a071fe04",
x"fe842783",
x"2783cf89",
x"8713fe44",
x"22230017",
x"17c1fee4",
x"071397a2",
x"8e2303a0",
x"2783fce7",
x"2703fe84",
x"97bafb84",
x"0007c783",
x"f7938391",
x"873e0ff7",
x"fec42783",
x"2783973e",
x"8693fe44",
x"22230017",
x"4703fed4",
x"17c10007",
x"8e2397a2",
x"2783fce7",
x"2703fe84",
x"97bafb84",
x"0007c783",
x"27038bbd",
x"973efec4",
x"fe442783",
x"00178693",
x"fed42223",
x"00074703",
x"97a217c1",
x"fce78e23",
x"fe842783",
x"24230785",
x"2703fef4",
x"4795fe84",
x"f6e7d8e3",
x"fac42783",
x"e7958bc1",
x"2783a819",
x"8713fbc4",
x"2e230017",
x"0713fae4",
x"80230200",
x"278300e7",
x"8713fb44",
x"2a23fff7",
x"2703fae4",
x"4ee3fe44",
x"2423fcf7",
x"a025fe04",
x"fbc42783",
x"00178713",
x"fae42e23",
x"fe842703",
x"97221741",
x"fdc74703",
x"00e78023",
x"fe842783",
x"24230785",
x"2703fef4",
x"2783fe84",
x"49e3fe44",
x"a819fcf7",
x"fbc42783",
x"00178713",
x"fae42e23",
x"02000713",
x"00e78023",
x"fb442783",
x"fff78713",
x"fae42a23",
x"fe442703",
x"fcf74ee3",
x"fbc42783",
x"4476853e",
x"80826125",
x"cea2711d",
x"2e231080",
x"2c23faa4",
x"2a23fab4",
x"2823fac4",
x"2623fad4",
x"2223fae4",
x"2623fe04",
x"a281fe04",
x"fec42783",
x"2783cf89",
x"8713fe44",
x"22230017",
x"17c1fee4",
x"071397a2",
x"8e2302e0",
x"2783fce7",
x"2703fec4",
x"97bafb84",
x"0007c783",
x"fef42423",
x"fe842783",
x"a703e385",
x"278380c1",
x"8693fe44",
x"22230017",
x"4703fed4",
x"17c10007",
x"8e2397a2",
x"a0cdfce7",
x"fe842703",
x"06300793",
x"06e7db63",
x"80c1a783",
x"fe842683",
x"06400713",
x"02e6c733",
x"2783973e",
x"8693fe44",
x"22230017",
x"4703fed4",
x"17c10007",
x"8e2397a2",
x"2703fce7",
x"0793fe84",
x"67b30640",
x"242302f7",
x"a783fef4",
x"268380c1",
x"4729fe84",
x"02e6c733",
x"2783973e",
x"8693fe44",
x"22230017",
x"4703fed4",
x"17c10007",
x"8e2397a2",
x"2703fce7",
x"47a9fe84",
x"02f767b3",
x"fef42423",
x"2703a089",
x"47a5fe84",
x"02e7dd63",
x"80c1a783",
x"fe842683",
x"c7334729",
x"973e02e6",
x"fe442783",
x"00178693",
x"fed42223",
x"00074703",
x"97a217c1",
x"fce78e23",
x"fe842703",
x"67b347a9",
x"242302f7",
x"a703fef4",
x"278380c1",
x"973efe84",
x"fe442783",
x"00178693",
x"fed42223",
x"00074703",
x"97a217c1",
x"fce78e23",
x"fec42783",
x"26230785",
x"2703fef4",
x"478dfec4",
x"eae7dee3",
x"fac42783",
x"e7958bc1",
x"2783a819",
x"8713fbc4",
x"2e230017",
x"0713fae4",
x"80230200",
x"278300e7",
x"8713fb44",
x"2a23fff7",
x"2703fae4",
x"4ee3fe44",
x"2623fcf7",
x"a025fe04",
x"fbc42783",
x"00178713",
x"fae42e23",
x"fec42703",
x"97221741",
x"fdc74703",
x"00e78023",
x"fec42783",
x"26230785",
x"2703fef4",
x"2783fec4",
x"49e3fe44",
x"a819fcf7",
x"fbc42783",
x"00178713",
x"fae42e23",
x"02000713",
x"00e78023",
x"fb442783",
x"fff78713",
x"fae42a23",
x"fe442703",
x"fcf74ee3",
x"fbc42783",
x"4476853e",
x"80826125",
x"c686715d",
x"0880c4a2",
x"faa42e23",
x"fab42c23",
x"fac42a23",
x"fbc42783",
x"fef42023",
x"2783a319",
x"c703fb84",
x"07930007",
x"0f630250",
x"270300f7",
x"2783fb84",
x"8693fe04",
x"20230017",
x"4703fed4",
x"80230007",
x"a9c900e7",
x"fc042c23",
x"fb842783",
x"2c230785",
x"2783faf4",
x"c783fb84",
x"17810007",
x"6d634741",
x"971304f7",
x"67a10027",
x"59878793",
x"439c97ba",
x"27838782",
x"e793fd84",
x"2c230107",
x"b7e9fcf4",
x"fd842783",
x"0047e793",
x"fcf42c23",
x"2783bf75",
x"e793fd84",
x"2c230087",
x"b77dfcf4",
x"fd842783",
x"0207e793",
x"fcf42c23",
x"2783b745",
x"e793fd84",
x"2c230017",
x"bf49fcf4",
x"2a2357fd",
x"2783fcf4",
x"c703fb84",
x"07930007",
x"f26302f0",
x"278302e7",
x"c703fb84",
x"07930007",
x"ea630390",
x"079300e7",
x"853efb84",
x"82fff0ef",
x"fca42a23",
x"2783a0b9",
x"c703fb84",
x"07930007",
x"106302a0",
x"278304f7",
x"0785fb84",
x"faf42c23",
x"fb442783",
x"00478713",
x"fae42a23",
x"2a23439c",
x"2783fcf4",
x"de63fd44",
x"27830007",
x"07b3fd44",
x"2a2340f0",
x"2783fcf4",
x"e793fd84",
x"2c230107",
x"57fdfcf4",
x"fcf42823",
x"fb842783",
x"0007c703",
x"02e00793",
x"06f71b63",
x"fb842783",
x"2c230785",
x"2783faf4",
x"c703fb84",
x"07930007",
x"f26302f0",
x"278302e7",
x"c703fb84",
x"07930007",
x"ea630390",
x"079300e7",
x"853efb84",
x"f92ff0ef",
x"fca42823",
x"2783a03d",
x"c703fb84",
x"07930007",
x"106302a0",
x"278302f7",
x"0785fb84",
x"faf42c23",
x"fb442783",
x"00478713",
x"fae42a23",
x"2823439c",
x"2783fcf4",
x"d463fd04",
x"28230007",
x"57fdfc04",
x"fcf42623",
x"fb842783",
x"0007c703",
x"06c00793",
x"00f70a63",
x"fb842783",
x"0007c703",
x"04c00793",
x"00f71d63",
x"fb842783",
x"0007c783",
x"fcf42623",
x"fb842783",
x"2c230785",
x"47a9faf4",
x"fef42223",
x"fb842783",
x"0007c783",
x"fbf78793",
x"03700713",
x"22f76e63",
x"00279713",
x"879367a1",
x"97ba5dc7",
x"8782439c",
x"fd842783",
x"e78d8bc1",
x"2783a819",
x"8713fe04",
x"20230017",
x"0713fee4",
x"80230200",
x"278300e7",
x"17fdfd44",
x"fcf42a23",
x"fd442783",
x"fcf04fe3",
x"fb442783",
x"00478713",
x"fae42a23",
x"27834394",
x"8713fe04",
x"20230017",
x"f713fee4",
x"80230ff6",
x"a81900e7",
x"fe042783",
x"00178713",
x"fee42023",
x"02000713",
x"00e78023",
x"fd442783",
x"2a2317fd",
x"2783fcf4",
x"4fe3fd44",
x"ac8dfcf0",
x"fb442783",
x"00478713",
x"fae42a23",
x"2e23439c",
x"2783fcf4",
x"e791fdc4",
x"879367a1",
x"2e235907",
x"2783fcf4",
x"85befd04",
x"fdc42503",
x"df4ff0ef",
x"242387aa",
x"2783fcf4",
x"8bc1fd84",
x"a819e795",
x"fe042783",
x"00178713",
x"fee42023",
x"02000713",
x"00e78023",
x"fd442783",
x"fff78713",
x"fce42a23",
x"fc842703",
x"fcf74ee3",
x"fe042423",
x"2703a035",
x"0793fdc4",
x"2e230017",
x"2783fcf4",
x"8693fe04",
x"20230017",
x"4703fed4",
x"80230007",
x"278300e7",
x"0785fe84",
x"fef42423",
x"fe842703",
x"fc842783",
x"fcf747e3",
x"2783a819",
x"8713fe04",
x"20230017",
x"0713fee4",
x"80230200",
x"278300e7",
x"8713fd44",
x"2a23fff7",
x"2703fce4",
x"4ee3fc84",
x"a24dfcf7",
x"fd442703",
x"1b6357fd",
x"47a100f7",
x"fcf42a23",
x"fd842783",
x"0017e793",
x"fcf42c23",
x"fb442783",
x"00478713",
x"fae42a23",
x"85be439c",
x"fd842783",
x"fd042703",
x"fd442683",
x"25034641",
x"f0effe04",
x"2023dccf",
x"aaa9fea4",
x"fd842783",
x"0407e793",
x"fcf42c23",
x"fcc42703",
x"06c00793",
x"02f71763",
x"fb442783",
x"00478713",
x"fae42a23",
x"2703439c",
x"2683fd84",
x"2603fd04",
x"85befd44",
x"fe042503",
x"88bff0ef",
x"fea42023",
x"2783aa21",
x"8713fb44",
x"2a230047",
x"439cfae4",
x"fd842703",
x"fd042683",
x"fd442603",
x"250385be",
x"3ac9fe04",
x"fea42023",
x"47a1a8c5",
x"fef42223",
x"2783a8ad",
x"e793fd84",
x"2c230407",
x"47c1fcf4",
x"fef42223",
x"2783a09d",
x"e793fd84",
x"2c230027",
x"a899fcf4",
x"fb842783",
x"0007c703",
x"02500793",
x"00f70c63",
x"fe042783",
x"00178713",
x"fee42023",
x"02500713",
x"00e78023",
x"fb842783",
x"0007c783",
x"2703cf91",
x"2783fb84",
x"8693fe04",
x"20230017",
x"4703fed4",
x"80230007",
x"a8bd00e7",
x"fb842783",
x"2c2317fd",
x"a88dfaf4",
x"27030001",
x"0793fcc4",
x"1c6306c0",
x"278300f7",
x"8713fb44",
x"2a230047",
x"439cfae4",
x"fef42623",
x"2783a805",
x"8b89fd84",
x"2783cb99",
x"8713fb44",
x"2a230047",
x"439cfae4",
x"fef42623",
x"2783a811",
x"8713fb44",
x"2a230047",
x"439cfae4",
x"fef42623",
x"fec42583",
x"fd842783",
x"fd042703",
x"fd442683",
x"fe442603",
x"fe042503",
x"c72ff0ef",
x"fea42023",
x"fb842783",
x"2c230785",
x"2783faf4",
x"c783fb84",
x"9ae30007",
x"2783ae07",
x"8023fe04",
x"27030007",
x"2783fe04",
x"07b3fbc4",
x"853e40f7",
x"442640b6",
x"80826161",
x"ce061101",
x"1000cc22",
x"07a387aa",
x"4703fef4",
x"47a9fef4",
x"00f71563",
x"c0ef4535",
x"4783bc5f",
x"853efef4",
x"bbbfc0ef",
x"40f20001",
x"61054462",
x"714d8082",
x"12112623",
x"12812423",
x"2e231a00",
x"c04ceca4",
x"c454c410",
x"c85cc818",
x"01042c23",
x"01142e23",
x"fe042423",
x"02040793",
x"ecf42c23",
x"ed842783",
x"22231791",
x"2703eef4",
x"0793ee44",
x"863aee84",
x"edc42583",
x"3c2d853e",
x"ee840793",
x"fef42623",
x"2783a00d",
x"c783fec4",
x"853e0007",
x"27833f85",
x"0785fe84",
x"fef42423",
x"fec42783",
x"26230785",
x"2783fef4",
x"c783fec4",
x"ffe10007",
x"fe842783",
x"2083853e",
x"240312c1",
x"61711281",
x"11018082",
x"cc22ce06",
x"26231000",
x"2423fea4",
x"2783feb4",
x"8793fec4",
x"25830427",
x"853efe84",
x"b89fe0ef",
x"40f20001",
x"61054462",
x"11018082",
x"cc22ce06",
x"26231000",
x"2783fea4",
x"8793fec4",
x"853e0427",
x"c1ffe0ef",
x"40f20001",
x"61054462",
x"711d8082",
x"cca2ce86",
x"45091080",
x"f00fc0ef",
x"fea42623",
x"f30fc0ef",
x"859367f1",
x"25032007",
x"c0effec4",
x"c0efa6df",
x"07938dbf",
x"2583fa44",
x"853efec4",
x"67a53fbd",
x"52a78793",
x"fef42423",
x"851367a1",
x"c0ef6bc7",
x"0713a6df",
x"2783fa44",
x"2583fe84",
x"853afec4",
x"07939782",
x"853efa44",
x"47813fbd",
x"40f6853e",
x"61254466",
x"00008082",
x"3340d4b0",
x"e7146a79",
x"0000e3c1",
x"1199be52",
x"1fd75608",
x"00000747",
x"39bf5e47",
x"8e3ae5a4",
x"00008d84",
x"00008420",
x"00008428",
x"00008430",
x"00008438",
x"00008440",
x"0000844c",
x"00008458",
x"00008464",
x"00008470",
x"0000847c",
x"00008488",
x"00008494",
x"000084a0",
x"000084ac",
x"000084b8",
x"000084c4",
x"00000000",
x"00000066",
x"0000000a",
x"00000001",
x"00008540",
x"00008568"
);
end neorv32_application_image;
